// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module conv2d_15_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h0001;
    tile_memory[  1] = 16'h2000;
    tile_memory[  2] = 16'h0202;
    tile_memory[  3] = 16'h00E0;
    tile_memory[  4] = 16'h8700;
    tile_memory[  5] = 16'h0006;
    tile_memory[  6] = 16'h1E04;
    tile_memory[  7] = 16'h0200;
    tile_memory[  8] = 16'h0F06;
    tile_memory[  9] = 16'h1F1F;
    tile_memory[ 10] = 16'h7070;
    tile_memory[ 11] = 16'h2165;
    tile_memory[ 12] = 16'h0480;
    tile_memory[ 13] = 16'h0686;
    tile_memory[ 14] = 16'h0E86;
    tile_memory[ 15] = 16'h040C;
    tile_memory[ 16] = 16'h7FFF;
    tile_memory[ 17] = 16'hEB3F;
    tile_memory[ 18] = 16'hEFFF;
    tile_memory[ 19] = 16'hBFA7;
    tile_memory[ 20] = 16'hFB78;
    tile_memory[ 21] = 16'h020F;
    tile_memory[ 22] = 16'hFF06;
    tile_memory[ 23] = 16'h07FF;
    tile_memory[ 24] = 16'h606C;
    tile_memory[ 25] = 16'h2121;
    tile_memory[ 26] = 16'h9C80;
    tile_memory[ 27] = 16'hC808;
    tile_memory[ 28] = 16'hC3C0;
    tile_memory[ 29] = 16'hE3A3;
    tile_memory[ 30] = 16'hC3D6;
    tile_memory[ 31] = 16'h8383;
    tile_memory[ 32] = 16'h0F4E;
    tile_memory[ 33] = 16'h4C46;
    tile_memory[ 34] = 16'hFC2C;
    tile_memory[ 35] = 16'h06FE;
    tile_memory[ 36] = 16'h8000;
    tile_memory[ 37] = 16'h0800;
    tile_memory[ 38] = 16'h0C04;
    tile_memory[ 39] = 16'h000C;
    tile_memory[ 40] = 16'hEF6F;
    tile_memory[ 41] = 16'h22FF;
    tile_memory[ 42] = 16'hF0E0;
    tile_memory[ 43] = 16'hF0F4;
    tile_memory[ 44] = 16'h3EB6;
    tile_memory[ 45] = 16'h040C;
    tile_memory[ 46] = 16'h6D00;
    tile_memory[ 47] = 16'hEDED;
    tile_memory[ 48] = 16'h1620;
    tile_memory[ 49] = 16'h4000;
    tile_memory[ 50] = 16'h0409;
    tile_memory[ 51] = 16'h0606;
    tile_memory[ 52] = 16'hC7DD;
    tile_memory[ 53] = 16'h1800;
    tile_memory[ 54] = 16'hA03C;
    tile_memory[ 55] = 16'h79F8;
    tile_memory[ 56] = 16'hD3C1;
    tile_memory[ 57] = 16'hF6F2;
    tile_memory[ 58] = 16'hC0F2;
    tile_memory[ 59] = 16'h8080;
    tile_memory[ 60] = 16'h0004;
    tile_memory[ 61] = 16'h0002;
    tile_memory[ 62] = 16'h1000;
    tile_memory[ 63] = 16'h000A;
    tile_memory[ 64] = 16'hFCF8;
    tile_memory[ 65] = 16'hE1E4;
    tile_memory[ 66] = 16'hCD63;
    tile_memory[ 67] = 16'hFD3D;
    tile_memory[ 68] = 16'h099F;
    tile_memory[ 69] = 16'hCB04;
    tile_memory[ 70] = 16'h9FB9;
    tile_memory[ 71] = 16'h70B6;
    tile_memory[ 72] = 16'h2F06;
    tile_memory[ 73] = 16'h8000;
    tile_memory[ 74] = 16'h20C4;
    tile_memory[ 75] = 16'hFF00;
    tile_memory[ 76] = 16'h1C00;
    tile_memory[ 77] = 16'h080C;
    tile_memory[ 78] = 16'h980C;
    tile_memory[ 79] = 16'h0C0E;
    tile_memory[ 80] = 16'h0706;
    tile_memory[ 81] = 16'hFE7F;
    tile_memory[ 82] = 16'hFE7E;
    tile_memory[ 83] = 16'hDE9E;
    tile_memory[ 84] = 16'h2000;
    tile_memory[ 85] = 16'h220F;
    tile_memory[ 86] = 16'hE600;
    tile_memory[ 87] = 16'hFBF9;
    tile_memory[ 88] = 16'hFFF8;
    tile_memory[ 89] = 16'h0A8C;
    tile_memory[ 90] = 16'hFDBE;
    tile_memory[ 91] = 16'h021F;
    tile_memory[ 92] = 16'hC3C5;
    tile_memory[ 93] = 16'h7836;
    tile_memory[ 94] = 16'h747C;
    tile_memory[ 95] = 16'h0060;
    tile_memory[ 96] = 16'h80E0;
    tile_memory[ 97] = 16'h0CA6;
    tile_memory[ 98] = 16'h9800;
    tile_memory[ 99] = 16'h0602;
    tile_memory[100] = 16'hE6E0;
    tile_memory[101] = 16'h2002;
    tile_memory[102] = 16'h6A78;
    tile_memory[103] = 16'h7F4E;
    tile_memory[104] = 16'hFF6F;
    tile_memory[105] = 16'h2EFF;
    tile_memory[106] = 16'hF5E0;
    tile_memory[107] = 16'h0008;
    tile_memory[108] = 16'hDFFF;
    tile_memory[109] = 16'h0006;
    tile_memory[110] = 16'h0800;
    tile_memory[111] = 16'h0101;
    tile_memory[112] = 16'h1660;
    tile_memory[113] = 16'h6000;
    tile_memory[114] = 16'h0804;
    tile_memory[115] = 16'h0010;
    tile_memory[116] = 16'h7900;
    tile_memory[117] = 16'hF878;
    tile_memory[118] = 16'hFCF0;
    tile_memory[119] = 16'h406C;
    tile_memory[120] = 16'h0F06;
    tile_memory[121] = 16'h1200;
    tile_memory[122] = 16'h0201;
    tile_memory[123] = 16'h0F38;
    tile_memory[124] = 16'hA200;
    tile_memory[125] = 16'h0002;
    tile_memory[126] = 16'h1300;
    tile_memory[127] = 16'h0003;
    tile_memory[128] = 16'h0F0C;
    tile_memory[129] = 16'h3F37;
    tile_memory[130] = 16'h073C;
    tile_memory[131] = 16'h8AEE;
    tile_memory[132] = 16'hFFFF;
    tile_memory[133] = 16'hFEFF;
    tile_memory[134] = 16'hD7FF;
    tile_memory[135] = 16'hFEF3;
    tile_memory[136] = 16'h1400;
    tile_memory[137] = 16'h0020;
    tile_memory[138] = 16'h0500;
    tile_memory[139] = 16'h4840;
    tile_memory[140] = 16'h0430;
    tile_memory[141] = 16'h0C00;
    tile_memory[142] = 16'h0400;
    tile_memory[143] = 16'h0004;
    tile_memory[144] = 16'h9F4F;
    tile_memory[145] = 16'hBFBF;
    tile_memory[146] = 16'hE7EC;
    tile_memory[147] = 16'hF7F7;
    tile_memory[148] = 16'h8000;
    tile_memory[149] = 16'h0307;
    tile_memory[150] = 16'hD404;
    tile_memory[151] = 16'h0383;
    tile_memory[152] = 16'hBF0F;
    tile_memory[153] = 16'h3FFF;
    tile_memory[154] = 16'hFCFE;
    tile_memory[155] = 16'h86E8;
    tile_memory[156] = 16'h2810;
    tile_memory[157] = 16'h8000;
    tile_memory[158] = 16'h6404;
    tile_memory[159] = 16'h7C1C;
    tile_memory[160] = 16'hDFFF;
    tile_memory[161] = 16'h8687;
    tile_memory[162] = 16'hC0C0;
    tile_memory[163] = 16'h4001;
    tile_memory[164] = 16'hF766;
    tile_memory[165] = 16'h00FF;
    tile_memory[166] = 16'hEEE1;
    tile_memory[167] = 16'h6FE0;
    tile_memory[168] = 16'h0804;
    tile_memory[169] = 16'h0707;
    tile_memory[170] = 16'h0177;
    tile_memory[171] = 16'h0606;
    tile_memory[172] = 16'h3820;
    tile_memory[173] = 16'h0020;
    tile_memory[174] = 16'h9C00;
    tile_memory[175] = 16'h001C;
    tile_memory[176] = 16'h7F4F;
    tile_memory[177] = 16'h7F7F;
    tile_memory[178] = 16'hE0E0;
    tile_memory[179] = 16'h0EFE;
    tile_memory[180] = 16'h3F4C;
    tile_memory[181] = 16'hFFFF;
    tile_memory[182] = 16'hF6FF;
    tile_memory[183] = 16'hF8F6;
    tile_memory[184] = 16'h0C0C;
    tile_memory[185] = 16'h3737;
    tile_memory[186] = 16'h0038;
    tile_memory[187] = 16'h0606;
    tile_memory[188] = 16'h001F;
    tile_memory[189] = 16'h0118;
    tile_memory[190] = 16'h4838;
    tile_memory[191] = 16'h1001;
    tile_memory[192] = 16'h1F0E;
    tile_memory[193] = 16'h233F;
    tile_memory[194] = 16'hE6FC;
    tile_memory[195] = 16'hE0F6;
    tile_memory[196] = 16'hFA70;
    tile_memory[197] = 16'hE8F0;
    tile_memory[198] = 16'h2240;
    tile_memory[199] = 16'h2900;
    tile_memory[200] = 16'h0202;
    tile_memory[201] = 16'h0002;
    tile_memory[202] = 16'h2000;
    tile_memory[203] = 16'h0068;
    tile_memory[204] = 16'h4F4F;
    tile_memory[205] = 16'h7F7F;
    tile_memory[206] = 16'hEC7E;
    tile_memory[207] = 16'hE9ED;
    tile_memory[208] = 16'h8200;
    tile_memory[209] = 16'h8404;
    tile_memory[210] = 16'h1000;
    tile_memory[211] = 16'h0280;
    tile_memory[212] = 16'hC1C7;
    tile_memory[213] = 16'hDFE7;
    tile_memory[214] = 16'hFFEB;
    tile_memory[215] = 16'hE1EC;
    tile_memory[216] = 16'h0A00;
    tile_memory[217] = 16'h2F3F;
    tile_memory[218] = 16'h165F;
    tile_memory[219] = 16'h0416;
    tile_memory[220] = 16'hFCED;
    tile_memory[221] = 16'hCDFC;
    tile_memory[222] = 16'h1F0F;
    tile_memory[223] = 16'hFFFF;
    tile_memory[224] = 16'hF670;
    tile_memory[225] = 16'hFCFC;
    tile_memory[226] = 16'hE7F1;
    tile_memory[227] = 16'h0026;
    tile_memory[228] = 16'h0006;
    tile_memory[229] = 16'h0C00;
    tile_memory[230] = 16'h1008;
    tile_memory[231] = 16'h0C00;
    tile_memory[232] = 16'hFF87;
    tile_memory[233] = 16'hFFFF;
    tile_memory[234] = 16'hFDE6;
    tile_memory[235] = 16'hF8F8;
    tile_memory[236] = 16'h0600;
    tile_memory[237] = 16'h00A0;
    tile_memory[238] = 16'h0C04;
    tile_memory[239] = 16'h0004;
    tile_memory[240] = 16'h0081;
    tile_memory[241] = 16'h2021;
    tile_memory[242] = 16'h0400;
    tile_memory[243] = 16'h0606;
    tile_memory[244] = 16'h1E50;
    tile_memory[245] = 16'h0100;
    tile_memory[246] = 16'hDF07;
    tile_memory[247] = 16'hFFFF;
    tile_memory[248] = 16'h0020;
    tile_memory[249] = 16'h0508;
    tile_memory[250] = 16'h0424;
    tile_memory[251] = 16'h0400;
    tile_memory[252] = 16'h1B08;
    tile_memory[253] = 16'hFE3F;
    tile_memory[254] = 16'hF6FE;
    tile_memory[255] = 16'h04E4;
  end

endmodule
