// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module fc_k_enc_1_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h0040;  // Neuron 0
    neuron_patterns[  1] = 16'h5981;  // Neuron 1
    neuron_patterns[  2] = 16'h0700;  // Neuron 2
    neuron_patterns[  3] = 16'h040D;  // Neuron 3
    neuron_patterns[  4] = 16'h5204;  // Neuron 4
    neuron_patterns[  5] = 16'h4080;  // Neuron 5
    neuron_patterns[  6] = 16'h0003;  // Neuron 6
    neuron_patterns[  7] = 16'h8804;  // Neuron 7
    neuron_patterns[  8] = 16'h0200;  // Neuron 8
    neuron_patterns[  9] = 16'h0340;  // Neuron 9
    neuron_patterns[ 10] = 16'h0000;  // Neuron 10
    neuron_patterns[ 11] = 16'h0000;  // Neuron 11
    neuron_patterns[ 12] = 16'h0380;  // Neuron 12
    neuron_patterns[ 13] = 16'h4120;  // Neuron 13
    neuron_patterns[ 14] = 16'h100C;  // Neuron 14
    neuron_patterns[ 15] = 16'h08E0;  // Neuron 15
    neuron_patterns[ 16] = 16'h0094;  // Neuron 16
    neuron_patterns[ 17] = 16'hC6A4;  // Neuron 17
    neuron_patterns[ 18] = 16'h0900;  // Neuron 18
    neuron_patterns[ 19] = 16'h0080;  // Neuron 19
    neuron_patterns[ 20] = 16'h0884;  // Neuron 20
    neuron_patterns[ 21] = 16'h0000;  // Neuron 21
    neuron_patterns[ 22] = 16'h0820;  // Neuron 22
    neuron_patterns[ 23] = 16'h8005;  // Neuron 23
    neuron_patterns[ 24] = 16'h4808;  // Neuron 24
    neuron_patterns[ 25] = 16'h0004;  // Neuron 25
    neuron_patterns[ 26] = 16'h1880;  // Neuron 26
    neuron_patterns[ 27] = 16'h4000;  // Neuron 27
    neuron_patterns[ 28] = 16'h0080;  // Neuron 28
    neuron_patterns[ 29] = 16'h0008;  // Neuron 29
    neuron_patterns[ 30] = 16'h8104;  // Neuron 30
    neuron_patterns[ 31] = 16'h0012;  // Neuron 31
    neuron_patterns[ 32] = 16'h0908;  // Neuron 32
    neuron_patterns[ 33] = 16'h6981;  // Neuron 33
    neuron_patterns[ 34] = 16'h0500;  // Neuron 34
    neuron_patterns[ 35] = 16'h0000;  // Neuron 35
    neuron_patterns[ 36] = 16'h78A4;  // Neuron 36
    neuron_patterns[ 37] = 16'h00A0;  // Neuron 37
    neuron_patterns[ 38] = 16'h0002;  // Neuron 38
    neuron_patterns[ 39] = 16'h4840;  // Neuron 39
    neuron_patterns[ 40] = 16'h4210;  // Neuron 40
    neuron_patterns[ 41] = 16'h0B40;  // Neuron 41
    neuron_patterns[ 42] = 16'h6000;  // Neuron 42
    neuron_patterns[ 43] = 16'h0600;  // Neuron 43
    neuron_patterns[ 44] = 16'h0380;  // Neuron 44
    neuron_patterns[ 45] = 16'h0020;  // Neuron 45
    neuron_patterns[ 46] = 16'h1008;  // Neuron 46
    neuron_patterns[ 47] = 16'h09E0;  // Neuron 47
    neuron_patterns[ 48] = 16'h0088;  // Neuron 48
    neuron_patterns[ 49] = 16'h040D;  // Neuron 49
    neuron_patterns[ 50] = 16'h0900;  // Neuron 50
    neuron_patterns[ 51] = 16'h0183;  // Neuron 51
    neuron_patterns[ 52] = 16'h08A0;  // Neuron 52
    neuron_patterns[ 53] = 16'h0800;  // Neuron 53
    neuron_patterns[ 54] = 16'h0920;  // Neuron 54
    neuron_patterns[ 55] = 16'h8005;  // Neuron 55
    neuron_patterns[ 56] = 16'h4000;  // Neuron 56
    neuron_patterns[ 57] = 16'h0000;  // Neuron 57
    neuron_patterns[ 58] = 16'h1801;  // Neuron 58
    neuron_patterns[ 59] = 16'h4200;  // Neuron 59
    neuron_patterns[ 60] = 16'h2080;  // Neuron 60
    neuron_patterns[ 61] = 16'h0108;  // Neuron 61
    neuron_patterns[ 62] = 16'hC100;  // Neuron 62
    neuron_patterns[ 63] = 16'h8012;  // Neuron 63
    neuron_patterns[ 64] = 16'h0941;  // Neuron 64
    neuron_patterns[ 65] = 16'h0080;  // Neuron 65
    neuron_patterns[ 66] = 16'h0000;  // Neuron 66
    neuron_patterns[ 67] = 16'h1001;  // Neuron 67
    neuron_patterns[ 68] = 16'h5804;  // Neuron 68
    neuron_patterns[ 69] = 16'h0020;  // Neuron 69
    neuron_patterns[ 70] = 16'h0000;  // Neuron 70
    neuron_patterns[ 71] = 16'h4800;  // Neuron 71
    neuron_patterns[ 72] = 16'h4311;  // Neuron 72
    neuron_patterns[ 73] = 16'h8141;  // Neuron 73
    neuron_patterns[ 74] = 16'h6100;  // Neuron 74
    neuron_patterns[ 75] = 16'h0480;  // Neuron 75
    neuron_patterns[ 76] = 16'h0380;  // Neuron 76
    neuron_patterns[ 77] = 16'h0020;  // Neuron 77
    neuron_patterns[ 78] = 16'h1008;  // Neuron 78
    neuron_patterns[ 79] = 16'h09E0;  // Neuron 79
    neuron_patterns[ 80] = 16'h0400;  // Neuron 80
    neuron_patterns[ 81] = 16'h800C;  // Neuron 81
    neuron_patterns[ 82] = 16'h0100;  // Neuron 82
    neuron_patterns[ 83] = 16'h4000;  // Neuron 83
    neuron_patterns[ 84] = 16'h0880;  // Neuron 84
    neuron_patterns[ 85] = 16'h0000;  // Neuron 85
    neuron_patterns[ 86] = 16'h0921;  // Neuron 86
    neuron_patterns[ 87] = 16'h8001;  // Neuron 87
    neuron_patterns[ 88] = 16'h0008;  // Neuron 88
    neuron_patterns[ 89] = 16'h0400;  // Neuron 89
    neuron_patterns[ 90] = 16'h0A80;  // Neuron 90
    neuron_patterns[ 91] = 16'h4000;  // Neuron 91
    neuron_patterns[ 92] = 16'h0080;  // Neuron 92
    neuron_patterns[ 93] = 16'h0308;  // Neuron 93
    neuron_patterns[ 94] = 16'h2080;  // Neuron 94
    neuron_patterns[ 95] = 16'h0032;  // Neuron 95
    neuron_patterns[ 96] = 16'h0901;  // Neuron 96
    neuron_patterns[ 97] = 16'hC184;  // Neuron 97
    neuron_patterns[ 98] = 16'h0000;  // Neuron 98
    neuron_patterns[ 99] = 16'h1400;  // Neuron 99
    neuron_patterns[100] = 16'h7804;  // Neuron 100
    neuron_patterns[101] = 16'h8411;  // Neuron 101
    neuron_patterns[102] = 16'h1000;  // Neuron 102
    neuron_patterns[103] = 16'h4904;  // Neuron 103
    neuron_patterns[104] = 16'h4000;  // Neuron 104
    neuron_patterns[105] = 16'hA441;  // Neuron 105
    neuron_patterns[106] = 16'h2100;  // Neuron 106
    neuron_patterns[107] = 16'h8040;  // Neuron 107
    neuron_patterns[108] = 16'h0A80;  // Neuron 108
    neuron_patterns[109] = 16'h0030;  // Neuron 109
    neuron_patterns[110] = 16'h0000;  // Neuron 110
    neuron_patterns[111] = 16'h08A0;  // Neuron 111
    neuron_patterns[112] = 16'h0221;  // Neuron 112
    neuron_patterns[113] = 16'h802D;  // Neuron 113
    neuron_patterns[114] = 16'h0100;  // Neuron 114
    neuron_patterns[115] = 16'h500A;  // Neuron 115
    neuron_patterns[116] = 16'h04A0;  // Neuron 116
    neuron_patterns[117] = 16'h0000;  // Neuron 117
    neuron_patterns[118] = 16'h0820;  // Neuron 118
    neuron_patterns[119] = 16'h0000;  // Neuron 119
    neuron_patterns[120] = 16'h0808;  // Neuron 120
    neuron_patterns[121] = 16'h0020;  // Neuron 121
    neuron_patterns[122] = 16'h48A0;  // Neuron 122
    neuron_patterns[123] = 16'h0880;  // Neuron 123
    neuron_patterns[124] = 16'h0000;  // Neuron 124
    neuron_patterns[125] = 16'h0248;  // Neuron 125
    neuron_patterns[126] = 16'h2084;  // Neuron 126
    neuron_patterns[127] = 16'h0020;  // Neuron 127
    neuron_patterns[128] = 16'h0940;  // Neuron 128
    neuron_patterns[129] = 16'hC184;  // Neuron 129
    neuron_patterns[130] = 16'h0420;  // Neuron 130
    neuron_patterns[131] = 16'h4400;  // Neuron 131
    neuron_patterns[132] = 16'h6B04;  // Neuron 132
    neuron_patterns[133] = 16'hC000;  // Neuron 133
    neuron_patterns[134] = 16'h00C2;  // Neuron 134
    neuron_patterns[135] = 16'h4B00;  // Neuron 135
    neuron_patterns[136] = 16'h8024;  // Neuron 136
    neuron_patterns[137] = 16'h2860;  // Neuron 137
    neuron_patterns[138] = 16'h0104;  // Neuron 138
    neuron_patterns[139] = 16'h8040;  // Neuron 139
    neuron_patterns[140] = 16'h1300;  // Neuron 140
    neuron_patterns[141] = 16'h0090;  // Neuron 141
    neuron_patterns[142] = 16'h1001;  // Neuron 142
    neuron_patterns[143] = 16'h0890;  // Neuron 143
    neuron_patterns[144] = 16'h22A9;  // Neuron 144
    neuron_patterns[145] = 16'h0024;  // Neuron 145
    neuron_patterns[146] = 16'h0900;  // Neuron 146
    neuron_patterns[147] = 16'h5009;  // Neuron 147
    neuron_patterns[148] = 16'h2060;  // Neuron 148
    neuron_patterns[149] = 16'h1808;  // Neuron 149
    neuron_patterns[150] = 16'hA821;  // Neuron 150
    neuron_patterns[151] = 16'h1800;  // Neuron 151
    neuron_patterns[152] = 16'h4808;  // Neuron 152
    neuron_patterns[153] = 16'h2021;  // Neuron 153
    neuron_patterns[154] = 16'h18C4;  // Neuron 154
    neuron_patterns[155] = 16'h4220;  // Neuron 155
    neuron_patterns[156] = 16'h1800;  // Neuron 156
    neuron_patterns[157] = 16'h4000;  // Neuron 157
    neuron_patterns[158] = 16'h0940;  // Neuron 158
    neuron_patterns[159] = 16'h0050;  // Neuron 159
    neuron_patterns[160] = 16'h1100;  // Neuron 160
    neuron_patterns[161] = 16'h4084;  // Neuron 161
    neuron_patterns[162] = 16'h0000;  // Neuron 162
    neuron_patterns[163] = 16'h0401;  // Neuron 163
    neuron_patterns[164] = 16'h480C;  // Neuron 164
    neuron_patterns[165] = 16'hC900;  // Neuron 165
    neuron_patterns[166] = 16'h0082;  // Neuron 166
    neuron_patterns[167] = 16'h4806;  // Neuron 167
    neuron_patterns[168] = 16'h9806;  // Neuron 168
    neuron_patterns[169] = 16'hA441;  // Neuron 169
    neuron_patterns[170] = 16'h0106;  // Neuron 170
    neuron_patterns[171] = 16'h1040;  // Neuron 171
    neuron_patterns[172] = 16'h1300;  // Neuron 172
    neuron_patterns[173] = 16'h0090;  // Neuron 173
    neuron_patterns[174] = 16'h0041;  // Neuron 174
    neuron_patterns[175] = 16'h0C10;  // Neuron 175
    neuron_patterns[176] = 16'h0388;  // Neuron 176
    neuron_patterns[177] = 16'h8E24;  // Neuron 177
    neuron_patterns[178] = 16'h0902;  // Neuron 178
    neuron_patterns[179] = 16'h5809;  // Neuron 179
    neuron_patterns[180] = 16'h0000;  // Neuron 180
    neuron_patterns[181] = 16'h0808;  // Neuron 181
    neuron_patterns[182] = 16'hCA11;  // Neuron 182
    neuron_patterns[183] = 16'h9000;  // Neuron 183
    neuron_patterns[184] = 16'h4C08;  // Neuron 184
    neuron_patterns[185] = 16'h2420;  // Neuron 185
    neuron_patterns[186] = 16'h9880;  // Neuron 186
    neuron_patterns[187] = 16'h4002;  // Neuron 187
    neuron_patterns[188] = 16'h1000;  // Neuron 188
    neuron_patterns[189] = 16'h0200;  // Neuron 189
    neuron_patterns[190] = 16'h2000;  // Neuron 190
    neuron_patterns[191] = 16'h8020;  // Neuron 191
    neuron_patterns[192] = 16'h1140;  // Neuron 192
    neuron_patterns[193] = 16'hC184;  // Neuron 193
    neuron_patterns[194] = 16'h0100;  // Neuron 194
    neuron_patterns[195] = 16'h0401;  // Neuron 195
    neuron_patterns[196] = 16'h728C;  // Neuron 196
    neuron_patterns[197] = 16'hC821;  // Neuron 197
    neuron_patterns[198] = 16'h0002;  // Neuron 198
    neuron_patterns[199] = 16'h0804;  // Neuron 199
    neuron_patterns[200] = 16'h5A00;  // Neuron 200
    neuron_patterns[201] = 16'h0441;  // Neuron 201
    neuron_patterns[202] = 16'h6104;  // Neuron 202
    neuron_patterns[203] = 16'h0080;  // Neuron 203
    neuron_patterns[204] = 16'h1380;  // Neuron 204
    neuron_patterns[205] = 16'h0080;  // Neuron 205
    neuron_patterns[206] = 16'h0000;  // Neuron 206
    neuron_patterns[207] = 16'h0840;  // Neuron 207
    neuron_patterns[208] = 16'h02D9;  // Neuron 208
    neuron_patterns[209] = 16'h8224;  // Neuron 209
    neuron_patterns[210] = 16'h0700;  // Neuron 210
    neuron_patterns[211] = 16'h5008;  // Neuron 211
    neuron_patterns[212] = 16'h0820;  // Neuron 212
    neuron_patterns[213] = 16'h0200;  // Neuron 213
    neuron_patterns[214] = 16'h0834;  // Neuron 214
    neuron_patterns[215] = 16'h9800;  // Neuron 215
    neuron_patterns[216] = 16'h0808;  // Neuron 216
    neuron_patterns[217] = 16'h0000;  // Neuron 217
    neuron_patterns[218] = 16'h1820;  // Neuron 218
    neuron_patterns[219] = 16'h4800;  // Neuron 219
    neuron_patterns[220] = 16'h0000;  // Neuron 220
    neuron_patterns[221] = 16'h4000;  // Neuron 221
    neuron_patterns[222] = 16'h0040;  // Neuron 222
    neuron_patterns[223] = 16'hA040;  // Neuron 223
    neuron_patterns[224] = 16'h1844;  // Neuron 224
    neuron_patterns[225] = 16'h6100;  // Neuron 225
    neuron_patterns[226] = 16'h0100;  // Neuron 226
    neuron_patterns[227] = 16'h0400;  // Neuron 227
    neuron_patterns[228] = 16'h7084;  // Neuron 228
    neuron_patterns[229] = 16'h8000;  // Neuron 229
    neuron_patterns[230] = 16'h0002;  // Neuron 230
    neuron_patterns[231] = 16'h4A00;  // Neuron 231
    neuron_patterns[232] = 16'h0000;  // Neuron 232
    neuron_patterns[233] = 16'h00C1;  // Neuron 233
    neuron_patterns[234] = 16'h6000;  // Neuron 234
    neuron_patterns[235] = 16'h0200;  // Neuron 235
    neuron_patterns[236] = 16'h1300;  // Neuron 236
    neuron_patterns[237] = 16'h4080;  // Neuron 237
    neuron_patterns[238] = 16'h0000;  // Neuron 238
    neuron_patterns[239] = 16'h08C1;  // Neuron 239
    neuron_patterns[240] = 16'h0050;  // Neuron 240
    neuron_patterns[241] = 16'h82A4;  // Neuron 241
    neuron_patterns[242] = 16'h0101;  // Neuron 242
    neuron_patterns[243] = 16'h0880;  // Neuron 243
    neuron_patterns[244] = 16'h0004;  // Neuron 244
    neuron_patterns[245] = 16'h0000;  // Neuron 245
    neuron_patterns[246] = 16'h0920;  // Neuron 246
    neuron_patterns[247] = 16'h8041;  // Neuron 247
    neuron_patterns[248] = 16'h4008;  // Neuron 248
    neuron_patterns[249] = 16'h2000;  // Neuron 249
    neuron_patterns[250] = 16'h1C00;  // Neuron 250
    neuron_patterns[251] = 16'h4800;  // Neuron 251
    neuron_patterns[252] = 16'h0000;  // Neuron 252
    neuron_patterns[253] = 16'h0008;  // Neuron 253
    neuron_patterns[254] = 16'h4000;  // Neuron 254
    neuron_patterns[255] = 16'h0030;  // Neuron 255
  end

endmodule
