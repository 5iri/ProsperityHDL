// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module attention_enc_0_kv_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'hEA62;
    tile_memory[  1] = 16'hDEDE;
    tile_memory[  2] = 16'h715F;
    tile_memory[  3] = 16'hF6F5;
    tile_memory[  4] = 16'h57D7;
    tile_memory[  5] = 16'h4747;
    tile_memory[  6] = 16'h97C7;
    tile_memory[  7] = 16'h1194;
    tile_memory[  8] = 16'h0511;
    tile_memory[  9] = 16'h9715;
    tile_memory[ 10] = 16'h9293;
    tile_memory[ 11] = 16'h9393;
    tile_memory[ 12] = 16'hC101;
    tile_memory[ 13] = 16'hEAE1;
    tile_memory[ 14] = 16'hCBEA;
    tile_memory[ 15] = 16'hC787;
    tile_memory[ 16] = 16'h44C6;
    tile_memory[ 17] = 16'h6F0D;
    tile_memory[ 18] = 16'hFEEB;
    tile_memory[ 19] = 16'hFE9C;
    tile_memory[ 20] = 16'h6E6E;
    tile_memory[ 21] = 16'h6C4C;
    tile_memory[ 22] = 16'hB12D;
    tile_memory[ 23] = 16'hB5B5;
    tile_memory[ 24] = 16'hA334;
    tile_memory[ 25] = 16'h87A7;
    tile_memory[ 26] = 16'h4CC4;
    tile_memory[ 27] = 16'h3A6A;
    tile_memory[ 28] = 16'h1D3E;
    tile_memory[ 29] = 16'hB115;
    tile_memory[ 30] = 16'hE9F9;
    tile_memory[ 31] = 16'h426B;
    tile_memory[ 32] = 16'hEA62;
    tile_memory[ 33] = 16'hDEDE;
    tile_memory[ 34] = 16'h71DF;
    tile_memory[ 35] = 16'hFEF5;
    tile_memory[ 36] = 16'h5FDF;
    tile_memory[ 37] = 16'h4747;
    tile_memory[ 38] = 16'h97C7;
    tile_memory[ 39] = 16'h199C;
    tile_memory[ 40] = 16'h0519;
    tile_memory[ 41] = 16'h9717;
    tile_memory[ 42] = 16'h9693;
    tile_memory[ 43] = 16'h9797;
    tile_memory[ 44] = 16'hC101;
    tile_memory[ 45] = 16'hEAE1;
    tile_memory[ 46] = 16'hCFEA;
    tile_memory[ 47] = 16'hC7C7;
    tile_memory[ 48] = 16'h44C6;
    tile_memory[ 49] = 16'h7F0D;
    tile_memory[ 50] = 16'hFEFB;
    tile_memory[ 51] = 16'hEF8D;
    tile_memory[ 52] = 16'h6F6F;
    tile_memory[ 53] = 16'h6C6D;
    tile_memory[ 54] = 16'hB12D;
    tile_memory[ 55] = 16'hB5B5;
    tile_memory[ 56] = 16'hE335;
    tile_memory[ 57] = 16'hC7E7;
    tile_memory[ 58] = 16'h4CC4;
    tile_memory[ 59] = 16'h3A6A;
    tile_memory[ 60] = 16'h3D3E;
    tile_memory[ 61] = 16'hF15D;
    tile_memory[ 62] = 16'hE9F9;
    tile_memory[ 63] = 16'h426B;
    tile_memory[ 64] = 16'hEAE2;
    tile_memory[ 65] = 16'hDEDE;
    tile_memory[ 66] = 16'hF1DF;
    tile_memory[ 67] = 16'hFEF7;
    tile_memory[ 68] = 16'h5FDF;
    tile_memory[ 69] = 16'h5757;
    tile_memory[ 70] = 16'hF7F7;
    tile_memory[ 71] = 16'h51F4;
    tile_memory[ 72] = 16'h0511;
    tile_memory[ 73] = 16'h9F1F;
    tile_memory[ 74] = 16'h969B;
    tile_memory[ 75] = 16'h9797;
    tile_memory[ 76] = 16'hC101;
    tile_memory[ 77] = 16'hEAE1;
    tile_memory[ 78] = 16'hCFEA;
    tile_memory[ 79] = 16'hCFC7;
    tile_memory[ 80] = 16'h4CCE;
    tile_memory[ 81] = 16'h7F0D;
    tile_memory[ 82] = 16'hFEFB;
    tile_memory[ 83] = 16'hEF8D;
    tile_memory[ 84] = 16'h6F6F;
    tile_memory[ 85] = 16'h6C6D;
    tile_memory[ 86] = 16'hB12D;
    tile_memory[ 87] = 16'hB5B5;
    tile_memory[ 88] = 16'hE335;
    tile_memory[ 89] = 16'hC7E7;
    tile_memory[ 90] = 16'h4CC4;
    tile_memory[ 91] = 16'h3A6A;
    tile_memory[ 92] = 16'h3D3E;
    tile_memory[ 93] = 16'hF15D;
    tile_memory[ 94] = 16'hE9F9;
    tile_memory[ 95] = 16'hC2EB;
    tile_memory[ 96] = 16'hFAFA;
    tile_memory[ 97] = 16'hDEDE;
    tile_memory[ 98] = 16'hF1DF;
    tile_memory[ 99] = 16'hFEF7;
    tile_memory[100] = 16'h5FDF;
    tile_memory[101] = 16'h5757;
    tile_memory[102] = 16'hB7F7;
    tile_memory[103] = 16'h19BC;
    tile_memory[104] = 16'h0519;
    tile_memory[105] = 16'h9F1F;
    tile_memory[106] = 16'h969F;
    tile_memory[107] = 16'hB797;
    tile_memory[108] = 16'hF121;
    tile_memory[109] = 16'hFBF1;
    tile_memory[110] = 16'hDFEA;
    tile_memory[111] = 16'hDFD7;
    tile_memory[112] = 16'h4ECE;
    tile_memory[113] = 16'h7F0F;
    tile_memory[114] = 16'hFEFB;
    tile_memory[115] = 16'hEF8D;
    tile_memory[116] = 16'h6F6F;
    tile_memory[117] = 16'h6D6D;
    tile_memory[118] = 16'hB12D;
    tile_memory[119] = 16'hB5B5;
    tile_memory[120] = 16'hF335;
    tile_memory[121] = 16'hC7F7;
    tile_memory[122] = 16'h4CC4;
    tile_memory[123] = 16'h3A6A;
    tile_memory[124] = 16'h3D3E;
    tile_memory[125] = 16'hF15D;
    tile_memory[126] = 16'hEBFB;
    tile_memory[127] = 16'hC6EF;
    tile_memory[128] = 16'hFAFA;
    tile_memory[129] = 16'hFEFE;
    tile_memory[130] = 16'h71FF;
    tile_memory[131] = 16'hFEF7;
    tile_memory[132] = 16'h5FDF;
    tile_memory[133] = 16'h5757;
    tile_memory[134] = 16'hFFFF;
    tile_memory[135] = 16'hD9FC;
    tile_memory[136] = 16'h0599;
    tile_memory[137] = 16'h9F1F;
    tile_memory[138] = 16'hD69F;
    tile_memory[139] = 16'hF7D7;
    tile_memory[140] = 16'hF1A1;
    tile_memory[141] = 16'hFBF1;
    tile_memory[142] = 16'hFFEA;
    tile_memory[143] = 16'hDFDF;
    tile_memory[144] = 16'h4ECE;
    tile_memory[145] = 16'h7F4F;
    tile_memory[146] = 16'hFEFB;
    tile_memory[147] = 16'hEF8D;
    tile_memory[148] = 16'h6F6F;
    tile_memory[149] = 16'h6D6D;
    tile_memory[150] = 16'hB32F;
    tile_memory[151] = 16'hB5B7;
    tile_memory[152] = 16'hF335;
    tile_memory[153] = 16'hC7F7;
    tile_memory[154] = 16'h5CD4;
    tile_memory[155] = 16'h3A7A;
    tile_memory[156] = 16'h3D3E;
    tile_memory[157] = 16'hF15D;
    tile_memory[158] = 16'hEFFF;
    tile_memory[159] = 16'hC6EF;
    tile_memory[160] = 16'hFAFA;
    tile_memory[161] = 16'hFEFE;
    tile_memory[162] = 16'h73FF;
    tile_memory[163] = 16'hFFF7;
    tile_memory[164] = 16'hDFDF;
    tile_memory[165] = 16'hC7D7;
    tile_memory[166] = 16'hFFEF;
    tile_memory[167] = 16'hD7FC;
    tile_memory[168] = 16'hD7D7;
    tile_memory[169] = 16'h9FDF;
    tile_memory[170] = 16'hD69F;
    tile_memory[171] = 16'hFFD7;
    tile_memory[172] = 16'hF9E9;
    tile_memory[173] = 16'hFBF9;
    tile_memory[174] = 16'hFFFA;
    tile_memory[175] = 16'hDFDF;
    tile_memory[176] = 16'hDEDE;
    tile_memory[177] = 16'hFF9F;
    tile_memory[178] = 16'hFEFB;
    tile_memory[179] = 16'hFF9F;
    tile_memory[180] = 16'hFF7F;
    tile_memory[181] = 16'hEDED;
    tile_memory[182] = 16'hFB6F;
    tile_memory[183] = 16'hF5FF;
    tile_memory[184] = 16'hF375;
    tile_memory[185] = 16'hCFFF;
    tile_memory[186] = 16'hDCDC;
    tile_memory[187] = 16'h7AFA;
    tile_memory[188] = 16'h3D3F;
    tile_memory[189] = 16'hF53D;
    tile_memory[190] = 16'hEFFF;
    tile_memory[191] = 16'hC6EF;
    tile_memory[192] = 16'hFBFA;
    tile_memory[193] = 16'hFFFF;
    tile_memory[194] = 16'h73FF;
    tile_memory[195] = 16'hFFF7;
    tile_memory[196] = 16'hDFDF;
    tile_memory[197] = 16'hC7D7;
    tile_memory[198] = 16'hFFEF;
    tile_memory[199] = 16'hD7FC;
    tile_memory[200] = 16'hD7D7;
    tile_memory[201] = 16'h9FDF;
    tile_memory[202] = 16'hD69F;
    tile_memory[203] = 16'hFFD7;
    tile_memory[204] = 16'hFFFD;
    tile_memory[205] = 16'hFFFF;
    tile_memory[206] = 16'hFFFE;
    tile_memory[207] = 16'hDFDF;
    tile_memory[208] = 16'hDEDE;
    tile_memory[209] = 16'hFFDF;
    tile_memory[210] = 16'hFEFF;
    tile_memory[211] = 16'hFF9D;
    tile_memory[212] = 16'hFF7F;
    tile_memory[213] = 16'hEDED;
    tile_memory[214] = 16'hFB6F;
    tile_memory[215] = 16'hF5FF;
    tile_memory[216] = 16'hF335;
    tile_memory[217] = 16'hEFFF;
    tile_memory[218] = 16'hDCFC;
    tile_memory[219] = 16'h7EFA;
    tile_memory[220] = 16'hBD3F;
    tile_memory[221] = 16'hF5FD;
    tile_memory[222] = 16'hEFFF;
    tile_memory[223] = 16'hC6EF;
    tile_memory[224] = 16'hFFBE;
    tile_memory[225] = 16'hFFFF;
    tile_memory[226] = 16'h7BFF;
    tile_memory[227] = 16'hFFF7;
    tile_memory[228] = 16'hDFDF;
    tile_memory[229] = 16'hE7F7;
    tile_memory[230] = 16'hFFEF;
    tile_memory[231] = 16'hFFFC;
    tile_memory[232] = 16'hD7DF;
    tile_memory[233] = 16'h9FDF;
    tile_memory[234] = 16'hD69F;
    tile_memory[235] = 16'hFFD7;
    tile_memory[236] = 16'hFFFD;
    tile_memory[237] = 16'hFFFF;
    tile_memory[238] = 16'hFFFE;
    tile_memory[239] = 16'hDFDF;
    tile_memory[240] = 16'hDEDE;
    tile_memory[241] = 16'hFF9F;
    tile_memory[242] = 16'hFFFF;
    tile_memory[243] = 16'hFF9F;
    tile_memory[244] = 16'hFF7F;
    tile_memory[245] = 16'hEFEF;
    tile_memory[246] = 16'hFB6F;
    tile_memory[247] = 16'hF5FF;
    tile_memory[248] = 16'hF3F5;
    tile_memory[249] = 16'hEFFF;
    tile_memory[250] = 16'hDEFE;
    tile_memory[251] = 16'h7EFA;
    tile_memory[252] = 16'hBD3F;
    tile_memory[253] = 16'hF7FF;
    tile_memory[254] = 16'hFFFF;
    tile_memory[255] = 16'hD6FF;
  end

endmodule
