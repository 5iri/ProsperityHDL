// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_v_enc_1_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h0220;
    tile_memory[  1] = 16'h29FC;
    tile_memory[  2] = 16'h56FB;
    tile_memory[  3] = 16'hAA29;
    tile_memory[  4] = 16'h0F9F;
    tile_memory[  5] = 16'h8B39;
    tile_memory[  6] = 16'h92D1;
    tile_memory[  7] = 16'hFDB4;
    tile_memory[  8] = 16'hA971;
    tile_memory[  9] = 16'hDBF5;
    tile_memory[ 10] = 16'h4077;
    tile_memory[ 11] = 16'hC9AB;
    tile_memory[ 12] = 16'h3BE7;
    tile_memory[ 13] = 16'hDB08;
    tile_memory[ 14] = 16'h6FC3;
    tile_memory[ 15] = 16'hB4E0;
    tile_memory[ 16] = 16'hFF02;
    tile_memory[ 17] = 16'h2335;
    tile_memory[ 18] = 16'hE294;
    tile_memory[ 19] = 16'h66F1;
    tile_memory[ 20] = 16'h1AA3;
    tile_memory[ 21] = 16'hD7D6;
    tile_memory[ 22] = 16'h4706;
    tile_memory[ 23] = 16'h3E2D;
    tile_memory[ 24] = 16'h485D;
    tile_memory[ 25] = 16'hCD40;
    tile_memory[ 26] = 16'h1C03;
    tile_memory[ 27] = 16'h09CB;
    tile_memory[ 28] = 16'h4D9B;
    tile_memory[ 29] = 16'h36AD;
    tile_memory[ 30] = 16'hA149;
    tile_memory[ 31] = 16'h213D;
    tile_memory[ 32] = 16'h60FA;
    tile_memory[ 33] = 16'h5459;
    tile_memory[ 34] = 16'h0954;
    tile_memory[ 35] = 16'hD20F;
    tile_memory[ 36] = 16'h41E8;
    tile_memory[ 37] = 16'hA724;
    tile_memory[ 38] = 16'h67C2;
    tile_memory[ 39] = 16'h6460;
    tile_memory[ 40] = 16'h38D2;
    tile_memory[ 41] = 16'hCAB8;
    tile_memory[ 42] = 16'hC983;
    tile_memory[ 43] = 16'hC409;
    tile_memory[ 44] = 16'hF940;
    tile_memory[ 45] = 16'h939C;
    tile_memory[ 46] = 16'h5B77;
    tile_memory[ 47] = 16'h8EB9;
    tile_memory[ 48] = 16'h0874;
    tile_memory[ 49] = 16'hB7E4;
    tile_memory[ 50] = 16'h6466;
    tile_memory[ 51] = 16'h6B0A;
    tile_memory[ 52] = 16'h130E;
    tile_memory[ 53] = 16'hC9D1;
    tile_memory[ 54] = 16'h91C3;
    tile_memory[ 55] = 16'hFD89;
    tile_memory[ 56] = 16'hC9CB;
    tile_memory[ 57] = 16'hC7E5;
    tile_memory[ 58] = 16'h2556;
    tile_memory[ 59] = 16'h6513;
    tile_memory[ 60] = 16'hAABB;
    tile_memory[ 61] = 16'h9388;
    tile_memory[ 62] = 16'hA049;
    tile_memory[ 63] = 16'h2546;
    tile_memory[ 64] = 16'hE604;
    tile_memory[ 65] = 16'h4643;
    tile_memory[ 66] = 16'hF9C3;
    tile_memory[ 67] = 16'h5420;
    tile_memory[ 68] = 16'h23A0;
    tile_memory[ 69] = 16'h5BDC;
    tile_memory[ 70] = 16'h670A;
    tile_memory[ 71] = 16'h04B3;
    tile_memory[ 72] = 16'h9EAC;
    tile_memory[ 73] = 16'hC511;
    tile_memory[ 74] = 16'h7E02;
    tile_memory[ 75] = 16'h317E;
    tile_memory[ 76] = 16'hD88B;
    tile_memory[ 77] = 16'h2839;
    tile_memory[ 78] = 16'h3B3A;
    tile_memory[ 79] = 16'hA88D;
    tile_memory[ 80] = 16'h6D32;
    tile_memory[ 81] = 16'hEF18;
    tile_memory[ 82] = 16'h6C96;
    tile_memory[ 83] = 16'hC315;
    tile_memory[ 84] = 16'h00A0;
    tile_memory[ 85] = 16'hF3B0;
    tile_memory[ 86] = 16'hACCF;
    tile_memory[ 87] = 16'hEF19;
    tile_memory[ 88] = 16'h0AAE;
    tile_memory[ 89] = 16'h9B2B;
    tile_memory[ 90] = 16'h9185;
    tile_memory[ 91] = 16'h223F;
    tile_memory[ 92] = 16'hD998;
    tile_memory[ 93] = 16'hEEBD;
    tile_memory[ 94] = 16'h5E3B;
    tile_memory[ 95] = 16'hCABD;
    tile_memory[ 96] = 16'hA2C2;
    tile_memory[ 97] = 16'h1BFE;
    tile_memory[ 98] = 16'h4E09;
    tile_memory[ 99] = 16'hEEBF;
    tile_memory[100] = 16'h396F;
    tile_memory[101] = 16'h8BB7;
    tile_memory[102] = 16'hF293;
    tile_memory[103] = 16'hD549;
    tile_memory[104] = 16'hEBF9;
    tile_memory[105] = 16'h93AF;
    tile_memory[106] = 16'hF873;
    tile_memory[107] = 16'h8D3B;
    tile_memory[108] = 16'h7B2F;
    tile_memory[109] = 16'hA28A;
    tile_memory[110] = 16'hED05;
    tile_memory[111] = 16'hB6D9;
    tile_memory[112] = 16'h578D;
    tile_memory[113] = 16'h64E3;
    tile_memory[114] = 16'h2BF0;
    tile_memory[115] = 16'h7736;
    tile_memory[116] = 16'h09F1;
    tile_memory[117] = 16'h06FC;
    tile_memory[118] = 16'hEEB6;
    tile_memory[119] = 16'hB16E;
    tile_memory[120] = 16'hA276;
    tile_memory[121] = 16'hCD55;
    tile_memory[122] = 16'hC400;
    tile_memory[123] = 16'h3850;
    tile_memory[124] = 16'hDBED;
    tile_memory[125] = 16'hEAE7;
    tile_memory[126] = 16'h07E1;
    tile_memory[127] = 16'h875D;
    tile_memory[128] = 16'hFD5E;
    tile_memory[129] = 16'hFE78;
    tile_memory[130] = 16'hBA4D;
    tile_memory[131] = 16'hD374;
    tile_memory[132] = 16'h77B3;
    tile_memory[133] = 16'hA926;
    tile_memory[134] = 16'hF0E7;
    tile_memory[135] = 16'hFED2;
    tile_memory[136] = 16'h4AAC;
    tile_memory[137] = 16'hDCFA;
    tile_memory[138] = 16'h2EC2;
    tile_memory[139] = 16'hF31F;
    tile_memory[140] = 16'hE98F;
    tile_memory[141] = 16'hD2FF;
    tile_memory[142] = 16'h717C;
    tile_memory[143] = 16'h8BE5;
    tile_memory[144] = 16'h25E0;
    tile_memory[145] = 16'hBD86;
    tile_memory[146] = 16'hDE39;
    tile_memory[147] = 16'h690A;
    tile_memory[148] = 16'h78C5;
    tile_memory[149] = 16'hABE4;
    tile_memory[150] = 16'hDDF7;
    tile_memory[151] = 16'hE7D2;
    tile_memory[152] = 16'hFF28;
    tile_memory[153] = 16'h8A1F;
    tile_memory[154] = 16'hD14E;
    tile_memory[155] = 16'h15A2;
    tile_memory[156] = 16'h3D75;
    tile_memory[157] = 16'hA04B;
    tile_memory[158] = 16'h4B79;
    tile_memory[159] = 16'h23DB;
    tile_memory[160] = 16'h3CF5;
    tile_memory[161] = 16'h21E5;
    tile_memory[162] = 16'h3194;
    tile_memory[163] = 16'h1D28;
    tile_memory[164] = 16'h6DE2;
    tile_memory[165] = 16'h757A;
    tile_memory[166] = 16'h7C69;
    tile_memory[167] = 16'hDBA5;
    tile_memory[168] = 16'h02E0;
    tile_memory[169] = 16'h5CDA;
    tile_memory[170] = 16'h4F03;
    tile_memory[171] = 16'hA26A;
    tile_memory[172] = 16'h6DAD;
    tile_memory[173] = 16'hB449;
    tile_memory[174] = 16'h2C36;
    tile_memory[175] = 16'h3B41;
    tile_memory[176] = 16'h5657;
    tile_memory[177] = 16'h9E92;
    tile_memory[178] = 16'h333F;
    tile_memory[179] = 16'h5766;
    tile_memory[180] = 16'hC908;
    tile_memory[181] = 16'hF7B2;
    tile_memory[182] = 16'hFD53;
    tile_memory[183] = 16'hDA4F;
    tile_memory[184] = 16'hD854;
    tile_memory[185] = 16'h1EE9;
    tile_memory[186] = 16'hF101;
    tile_memory[187] = 16'h8B49;
    tile_memory[188] = 16'hFDED;
    tile_memory[189] = 16'h13DC;
    tile_memory[190] = 16'h39D0;
    tile_memory[191] = 16'h6BAC;
    tile_memory[192] = 16'hE88B;
    tile_memory[193] = 16'h88C9;
    tile_memory[194] = 16'h0ECC;
    tile_memory[195] = 16'h89E4;
    tile_memory[196] = 16'hFECF;
    tile_memory[197] = 16'h6972;
    tile_memory[198] = 16'h795D;
    tile_memory[199] = 16'h478A;
    tile_memory[200] = 16'h1B3E;
    tile_memory[201] = 16'hF2ED;
    tile_memory[202] = 16'hA95F;
    tile_memory[203] = 16'hAA16;
    tile_memory[204] = 16'h356F;
    tile_memory[205] = 16'hD6BA;
    tile_memory[206] = 16'h1AB3;
    tile_memory[207] = 16'hE8E3;
    tile_memory[208] = 16'hEE54;
    tile_memory[209] = 16'h2C89;
    tile_memory[210] = 16'hA3E9;
    tile_memory[211] = 16'h0BA9;
    tile_memory[212] = 16'h8BBC;
    tile_memory[213] = 16'h6BFC;
    tile_memory[214] = 16'h473C;
    tile_memory[215] = 16'h09B3;
    tile_memory[216] = 16'h3079;
    tile_memory[217] = 16'hA704;
    tile_memory[218] = 16'h78E1;
    tile_memory[219] = 16'hEB78;
    tile_memory[220] = 16'h083D;
    tile_memory[221] = 16'h7851;
    tile_memory[222] = 16'h9C18;
    tile_memory[223] = 16'h64B7;
    tile_memory[224] = 16'h4EF0;
    tile_memory[225] = 16'hEB1F;
    tile_memory[226] = 16'h95EA;
    tile_memory[227] = 16'h2E4F;
    tile_memory[228] = 16'h3D57;
    tile_memory[229] = 16'hFB73;
    tile_memory[230] = 16'hF4C0;
    tile_memory[231] = 16'h6758;
    tile_memory[232] = 16'h6CF0;
    tile_memory[233] = 16'h2834;
    tile_memory[234] = 16'hE7E1;
    tile_memory[235] = 16'h569F;
    tile_memory[236] = 16'hA418;
    tile_memory[237] = 16'h1AEC;
    tile_memory[238] = 16'h5DC1;
    tile_memory[239] = 16'hCA53;
    tile_memory[240] = 16'h1240;
    tile_memory[241] = 16'h01CC;
    tile_memory[242] = 16'hDE3D;
    tile_memory[243] = 16'h8E1E;
    tile_memory[244] = 16'h3124;
    tile_memory[245] = 16'h4B7B;
    tile_memory[246] = 16'hB083;
    tile_memory[247] = 16'h4710;
    tile_memory[248] = 16'hE5A7;
    tile_memory[249] = 16'hBBA7;
    tile_memory[250] = 16'h2855;
    tile_memory[251] = 16'h4C1B;
    tile_memory[252] = 16'h39A7;
    tile_memory[253] = 16'hB89D;
    tile_memory[254] = 16'hCC8D;
    tile_memory[255] = 16'h3741;
  end

endmodule
