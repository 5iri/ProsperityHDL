// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module attention_enc_1_kv_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h0505;  // Neuron 0
    neuron_patterns[  1] = 16'h6624;  // Neuron 1
    neuron_patterns[  2] = 16'h4363;  // Neuron 2
    neuron_patterns[  3] = 16'hA421;  // Neuron 3
    neuron_patterns[  4] = 16'hCCE4;  // Neuron 4
    neuron_patterns[  5] = 16'h7FCF;  // Neuron 5
    neuron_patterns[  6] = 16'h3677;  // Neuron 6
    neuron_patterns[  7] = 16'h482C;  // Neuron 7
    neuron_patterns[  8] = 16'hD0D8;  // Neuron 8
    neuron_patterns[  9] = 16'h1A9A;  // Neuron 9
    neuron_patterns[ 10] = 16'h131B;  // Neuron 10
    neuron_patterns[ 11] = 16'h7515;  // Neuron 11
    neuron_patterns[ 12] = 16'hEAE7;  // Neuron 12
    neuron_patterns[ 13] = 16'h0F8F;  // Neuron 13
    neuron_patterns[ 14] = 16'hA7A7;  // Neuron 14
    neuron_patterns[ 15] = 16'h5FBD;  // Neuron 15
    neuron_patterns[ 16] = 16'hDB5B;  // Neuron 16
    neuron_patterns[ 17] = 16'h889A;  // Neuron 17
    neuron_patterns[ 18] = 16'h7070;  // Neuron 18
    neuron_patterns[ 19] = 16'h0270;  // Neuron 19
    neuron_patterns[ 20] = 16'hFA2A;  // Neuron 20
    neuron_patterns[ 21] = 16'hF0F8;  // Neuron 21
    neuron_patterns[ 22] = 16'h5A3A;  // Neuron 22
    neuron_patterns[ 23] = 16'hD3DA;  // Neuron 23
    neuron_patterns[ 24] = 16'hCFDD;  // Neuron 24
    neuron_patterns[ 25] = 16'h92DF;  // Neuron 25
    neuron_patterns[ 26] = 16'h4F93;  // Neuron 26
    neuron_patterns[ 27] = 16'h5F5F;  // Neuron 27
    neuron_patterns[ 28] = 16'h5353;  // Neuron 28
    neuron_patterns[ 29] = 16'hD5D3;  // Neuron 29
    neuron_patterns[ 30] = 16'hF5F5;  // Neuron 30
    neuron_patterns[ 31] = 16'h01B5;  // Neuron 31
    neuron_patterns[ 32] = 16'h8585;  // Neuron 32
    neuron_patterns[ 33] = 16'h6724;  // Neuron 33
    neuron_patterns[ 34] = 16'h4363;  // Neuron 34
    neuron_patterns[ 35] = 16'hF571;  // Neuron 35
    neuron_patterns[ 36] = 16'hCDF5;  // Neuron 36
    neuron_patterns[ 37] = 16'h7FCF;  // Neuron 37
    neuron_patterns[ 38] = 16'h3677;  // Neuron 38
    neuron_patterns[ 39] = 16'hC8A8;  // Neuron 39
    neuron_patterns[ 40] = 16'hD1D8;  // Neuron 40
    neuron_patterns[ 41] = 16'hDBDB;  // Neuron 41
    neuron_patterns[ 42] = 16'h93DB;  // Neuron 42
    neuron_patterns[ 43] = 16'hF595;  // Neuron 43
    neuron_patterns[ 44] = 16'hEAE7;  // Neuron 44
    neuron_patterns[ 45] = 16'h2FAF;  // Neuron 45
    neuron_patterns[ 46] = 16'hA6A7;  // Neuron 46
    neuron_patterns[ 47] = 16'h7DBC;  // Neuron 47
    neuron_patterns[ 48] = 16'hDB7B;  // Neuron 48
    neuron_patterns[ 49] = 16'h8C9A;  // Neuron 49
    neuron_patterns[ 50] = 16'h7C7C;  // Neuron 50
    neuron_patterns[ 51] = 16'h0378;  // Neuron 51
    neuron_patterns[ 52] = 16'hBB2B;  // Neuron 52
    neuron_patterns[ 53] = 16'hB0B8;  // Neuron 53
    neuron_patterns[ 54] = 16'hDB9B;  // Neuron 54
    neuron_patterns[ 55] = 16'hF3DB;  // Neuron 55
    neuron_patterns[ 56] = 16'hEFFD;  // Neuron 56
    neuron_patterns[ 57] = 16'hF2FF;  // Neuron 57
    neuron_patterns[ 58] = 16'h4FB3;  // Neuron 58
    neuron_patterns[ 59] = 16'h5D5D;  // Neuron 59
    neuron_patterns[ 60] = 16'h4353;  // Neuron 60
    neuron_patterns[ 61] = 16'hC7C7;  // Neuron 61
    neuron_patterns[ 62] = 16'h7FFF;  // Neuron 62
    neuron_patterns[ 63] = 16'h013D;  // Neuron 63
    neuron_patterns[ 64] = 16'h8585;  // Neuron 64
    neuron_patterns[ 65] = 16'h6724;  // Neuron 65
    neuron_patterns[ 66] = 16'hC3E3;  // Neuron 66
    neuron_patterns[ 67] = 16'hF7F1;  // Neuron 67
    neuron_patterns[ 68] = 16'hCFF7;  // Neuron 68
    neuron_patterns[ 69] = 16'h7FCF;  // Neuron 69
    neuron_patterns[ 70] = 16'hBE77;  // Neuron 70
    neuron_patterns[ 71] = 16'hE8AA;  // Neuron 71
    neuron_patterns[ 72] = 16'hF1D8;  // Neuron 72
    neuron_patterns[ 73] = 16'hFBFB;  // Neuron 73
    neuron_patterns[ 74] = 16'hB3FB;  // Neuron 74
    neuron_patterns[ 75] = 16'hF5B5;  // Neuron 75
    neuron_patterns[ 76] = 16'hEAE7;  // Neuron 76
    neuron_patterns[ 77] = 16'h2FAF;  // Neuron 77
    neuron_patterns[ 78] = 16'hA6A7;  // Neuron 78
    neuron_patterns[ 79] = 16'h7FBC;  // Neuron 79
    neuron_patterns[ 80] = 16'hDB7B;  // Neuron 80
    neuron_patterns[ 81] = 16'hC8DA;  // Neuron 81
    neuron_patterns[ 82] = 16'hF878;  // Neuron 82
    neuron_patterns[ 83] = 16'h8BF8;  // Neuron 83
    neuron_patterns[ 84] = 16'hFB3B;  // Neuron 84
    neuron_patterns[ 85] = 16'hF0F8;  // Neuron 85
    neuron_patterns[ 86] = 16'hDB9B;  // Neuron 86
    neuron_patterns[ 87] = 16'hF3DB;  // Neuron 87
    neuron_patterns[ 88] = 16'hEFFD;  // Neuron 88
    neuron_patterns[ 89] = 16'hF2FF;  // Neuron 89
    neuron_patterns[ 90] = 16'h4FB3;  // Neuron 90
    neuron_patterns[ 91] = 16'hDF5F;  // Neuron 91
    neuron_patterns[ 92] = 16'hC3D3;  // Neuron 92
    neuron_patterns[ 93] = 16'hC7C7;  // Neuron 93
    neuron_patterns[ 94] = 16'hFFFF;  // Neuron 94
    neuron_patterns[ 95] = 16'h01BD;  // Neuron 95
    neuron_patterns[ 96] = 16'h8787;  // Neuron 96
    neuron_patterns[ 97] = 16'h67A6;  // Neuron 97
    neuron_patterns[ 98] = 16'hC3E3;  // Neuron 98
    neuron_patterns[ 99] = 16'hF7F1;  // Neuron 99
    neuron_patterns[100] = 16'hEFF7;  // Neuron 100
    neuron_patterns[101] = 16'h7FEF;  // Neuron 101
    neuron_patterns[102] = 16'hBE77;  // Neuron 102
    neuron_patterns[103] = 16'hE9AA;  // Neuron 103
    neuron_patterns[104] = 16'hF9D9;  // Neuron 104
    neuron_patterns[105] = 16'hFBFB;  // Neuron 105
    neuron_patterns[106] = 16'hB3FB;  // Neuron 106
    neuron_patterns[107] = 16'hD5B5;  // Neuron 107
    neuron_patterns[108] = 16'hEAC7;  // Neuron 108
    neuron_patterns[109] = 16'hAFAF;  // Neuron 109
    neuron_patterns[110] = 16'hA6A7;  // Neuron 110
    neuron_patterns[111] = 16'h7FBC;  // Neuron 111
    neuron_patterns[112] = 16'hDF7F;  // Neuron 112
    neuron_patterns[113] = 16'hCCDA;  // Neuron 113
    neuron_patterns[114] = 16'hFC7C;  // Neuron 114
    neuron_patterns[115] = 16'h8BF8;  // Neuron 115
    neuron_patterns[116] = 16'hFB3B;  // Neuron 116
    neuron_patterns[117] = 16'hF2FA;  // Neuron 117
    neuron_patterns[118] = 16'hDB9B;  // Neuron 118
    neuron_patterns[119] = 16'hF3DB;  // Neuron 119
    neuron_patterns[120] = 16'hFFFD;  // Neuron 120
    neuron_patterns[121] = 16'hF6FF;  // Neuron 121
    neuron_patterns[122] = 16'h4FB7;  // Neuron 122
    neuron_patterns[123] = 16'hDF5F;  // Neuron 123
    neuron_patterns[124] = 16'hFBD3;  // Neuron 124
    neuron_patterns[125] = 16'hBFFF;  // Neuron 125
    neuron_patterns[126] = 16'h3FBF;  // Neuron 126
    neuron_patterns[127] = 16'h013D;  // Neuron 127
    neuron_patterns[128] = 16'h8787;  // Neuron 128
    neuron_patterns[129] = 16'h6766;  // Neuron 129
    neuron_patterns[130] = 16'hC3E3;  // Neuron 130
    neuron_patterns[131] = 16'hFDF9;  // Neuron 131
    neuron_patterns[132] = 16'hEDFD;  // Neuron 132
    neuron_patterns[133] = 16'h7FFF;  // Neuron 133
    neuron_patterns[134] = 16'h3E77;  // Neuron 134
    neuron_patterns[135] = 16'hE8AE;  // Neuron 135
    neuron_patterns[136] = 16'hF9D8;  // Neuron 136
    neuron_patterns[137] = 16'hFBFB;  // Neuron 137
    neuron_patterns[138] = 16'hB3FB;  // Neuron 138
    neuron_patterns[139] = 16'hF5B5;  // Neuron 139
    neuron_patterns[140] = 16'hEAE7;  // Neuron 140
    neuron_patterns[141] = 16'hAFAF;  // Neuron 141
    neuron_patterns[142] = 16'hA7A7;  // Neuron 142
    neuron_patterns[143] = 16'h7FBC;  // Neuron 143
    neuron_patterns[144] = 16'hDB7B;  // Neuron 144
    neuron_patterns[145] = 16'hDCDA;  // Neuron 145
    neuron_patterns[146] = 16'hFE7E;  // Neuron 146
    neuron_patterns[147] = 16'hCFFA;  // Neuron 147
    neuron_patterns[148] = 16'hFF3F;  // Neuron 148
    neuron_patterns[149] = 16'hF2FA;  // Neuron 149
    neuron_patterns[150] = 16'hDB9B;  // Neuron 150
    neuron_patterns[151] = 16'hF7DF;  // Neuron 151
    neuron_patterns[152] = 16'hEFFD;  // Neuron 152
    neuron_patterns[153] = 16'hF6FF;  // Neuron 153
    neuron_patterns[154] = 16'h4FF7;  // Neuron 154
    neuron_patterns[155] = 16'hDD5D;  // Neuron 155
    neuron_patterns[156] = 16'hFBDB;  // Neuron 156
    neuron_patterns[157] = 16'hB7FF;  // Neuron 157
    neuron_patterns[158] = 16'hBFBF;  // Neuron 158
    neuron_patterns[159] = 16'h01BD;  // Neuron 159
    neuron_patterns[160] = 16'hD797;  // Neuron 160
    neuron_patterns[161] = 16'h67E6;  // Neuron 161
    neuron_patterns[162] = 16'hC3E3;  // Neuron 162
    neuron_patterns[163] = 16'hFFF9;  // Neuron 163
    neuron_patterns[164] = 16'hEFFF;  // Neuron 164
    neuron_patterns[165] = 16'h7FFF;  // Neuron 165
    neuron_patterns[166] = 16'hBE77;  // Neuron 166
    neuron_patterns[167] = 16'hE9AA;  // Neuron 167
    neuron_patterns[168] = 16'hD9D9;  // Neuron 168
    neuron_patterns[169] = 16'hDBDB;  // Neuron 169
    neuron_patterns[170] = 16'hBBFB;  // Neuron 170
    neuron_patterns[171] = 16'hF5BD;  // Neuron 171
    neuron_patterns[172] = 16'hEEE7;  // Neuron 172
    neuron_patterns[173] = 16'hAFAF;  // Neuron 173
    neuron_patterns[174] = 16'hA7A7;  // Neuron 174
    neuron_patterns[175] = 16'h7FBC;  // Neuron 175
    neuron_patterns[176] = 16'hDF7B;  // Neuron 176
    neuron_patterns[177] = 16'hDDDF;  // Neuron 177
    neuron_patterns[178] = 16'hFF7F;  // Neuron 178
    neuron_patterns[179] = 16'h8FFB;  // Neuron 179
    neuron_patterns[180] = 16'hFF3F;  // Neuron 180
    neuron_patterns[181] = 16'hF2FE;  // Neuron 181
    neuron_patterns[182] = 16'hDB9B;  // Neuron 182
    neuron_patterns[183] = 16'hF7DF;  // Neuron 183
    neuron_patterns[184] = 16'hFFFD;  // Neuron 184
    neuron_patterns[185] = 16'hF6FF;  // Neuron 185
    neuron_patterns[186] = 16'hCFB7;  // Neuron 186
    neuron_patterns[187] = 16'hDFDF;  // Neuron 187
    neuron_patterns[188] = 16'hFBDB;  // Neuron 188
    neuron_patterns[189] = 16'hFFFF;  // Neuron 189
    neuron_patterns[190] = 16'hFFFF;  // Neuron 190
    neuron_patterns[191] = 16'h01FD;  // Neuron 191
    neuron_patterns[192] = 16'hC787;  // Neuron 192
    neuron_patterns[193] = 16'h67E6;  // Neuron 193
    neuron_patterns[194] = 16'hDBEB;  // Neuron 194
    neuron_patterns[195] = 16'hFDF9;  // Neuron 195
    neuron_patterns[196] = 16'hEDFD;  // Neuron 196
    neuron_patterns[197] = 16'h7FFF;  // Neuron 197
    neuron_patterns[198] = 16'h3E77;  // Neuron 198
    neuron_patterns[199] = 16'hEDAA;  // Neuron 199
    neuron_patterns[200] = 16'hFFDD;  // Neuron 200
    neuron_patterns[201] = 16'hFBFB;  // Neuron 201
    neuron_patterns[202] = 16'hBFFB;  // Neuron 202
    neuron_patterns[203] = 16'hF5BD;  // Neuron 203
    neuron_patterns[204] = 16'hEEE7;  // Neuron 204
    neuron_patterns[205] = 16'hAFAF;  // Neuron 205
    neuron_patterns[206] = 16'hA7A7;  // Neuron 206
    neuron_patterns[207] = 16'h7FBE;  // Neuron 207
    neuron_patterns[208] = 16'hDF7B;  // Neuron 208
    neuron_patterns[209] = 16'hDDDF;  // Neuron 209
    neuron_patterns[210] = 16'hFF7F;  // Neuron 210
    neuron_patterns[211] = 16'hCFFB;  // Neuron 211
    neuron_patterns[212] = 16'hFF3F;  // Neuron 212
    neuron_patterns[213] = 16'hF6FE;  // Neuron 213
    neuron_patterns[214] = 16'hDF9F;  // Neuron 214
    neuron_patterns[215] = 16'hF7DF;  // Neuron 215
    neuron_patterns[216] = 16'hEFFD;  // Neuron 216
    neuron_patterns[217] = 16'hF2FF;  // Neuron 217
    neuron_patterns[218] = 16'hDFB3;  // Neuron 218
    neuron_patterns[219] = 16'hDFDF;  // Neuron 219
    neuron_patterns[220] = 16'hFBDB;  // Neuron 220
    neuron_patterns[221] = 16'hFFFF;  // Neuron 221
    neuron_patterns[222] = 16'hFFFF;  // Neuron 222
    neuron_patterns[223] = 16'h01FF;  // Neuron 223
    neuron_patterns[224] = 16'h8787;  // Neuron 224
    neuron_patterns[225] = 16'h6FEF;  // Neuron 225
    neuron_patterns[226] = 16'hDBEB;  // Neuron 226
    neuron_patterns[227] = 16'hFFF9;  // Neuron 227
    neuron_patterns[228] = 16'hEFFF;  // Neuron 228
    neuron_patterns[229] = 16'h7FFF;  // Neuron 229
    neuron_patterns[230] = 16'hBE77;  // Neuron 230
    neuron_patterns[231] = 16'hEDAA;  // Neuron 231
    neuron_patterns[232] = 16'hFFDD;  // Neuron 232
    neuron_patterns[233] = 16'hFBFB;  // Neuron 233
    neuron_patterns[234] = 16'hBFFB;  // Neuron 234
    neuron_patterns[235] = 16'hF7BF;  // Neuron 235
    neuron_patterns[236] = 16'hEFFF;  // Neuron 236
    neuron_patterns[237] = 16'hAFAF;  // Neuron 237
    neuron_patterns[238] = 16'hB7B7;  // Neuron 238
    neuron_patterns[239] = 16'h7FBE;  // Neuron 239
    neuron_patterns[240] = 16'hFF7F;  // Neuron 240
    neuron_patterns[241] = 16'hCDDF;  // Neuron 241
    neuron_patterns[242] = 16'hFB7B;  // Neuron 242
    neuron_patterns[243] = 16'hCFFB;  // Neuron 243
    neuron_patterns[244] = 16'hFF3F;  // Neuron 244
    neuron_patterns[245] = 16'hF6FE;  // Neuron 245
    neuron_patterns[246] = 16'hDFBF;  // Neuron 246
    neuron_patterns[247] = 16'hF7DF;  // Neuron 247
    neuron_patterns[248] = 16'hFFFD;  // Neuron 248
    neuron_patterns[249] = 16'hF3FF;  // Neuron 249
    neuron_patterns[250] = 16'hCFF3;  // Neuron 250
    neuron_patterns[251] = 16'hDDDD;  // Neuron 251
    neuron_patterns[252] = 16'hFBDB;  // Neuron 252
    neuron_patterns[253] = 16'hFFFF;  // Neuron 253
    neuron_patterns[254] = 16'hFFFF;  // Neuron 254
    neuron_patterns[255] = 16'h01FF;  // Neuron 255
  end

endmodule
