// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module conv2d_0_sps_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'hFFFF;  // Neuron 0
    neuron_patterns[  1] = 16'hFFFF;  // Neuron 1
    neuron_patterns[  2] = 16'hFFFF;  // Neuron 2
    neuron_patterns[  3] = 16'hFFFF;  // Neuron 3
    neuron_patterns[  4] = 16'hFFFF;  // Neuron 4
    neuron_patterns[  5] = 16'hFFFF;  // Neuron 5
    neuron_patterns[  6] = 16'hFFFF;  // Neuron 6
    neuron_patterns[  7] = 16'hFFFF;  // Neuron 7
    neuron_patterns[  8] = 16'hFFFF;  // Neuron 8
    neuron_patterns[  9] = 16'hFFFF;  // Neuron 9
    neuron_patterns[ 10] = 16'hFFFF;  // Neuron 10
    neuron_patterns[ 11] = 16'hFFFF;  // Neuron 11
    neuron_patterns[ 12] = 16'hFFFF;  // Neuron 12
    neuron_patterns[ 13] = 16'hFFFF;  // Neuron 13
    neuron_patterns[ 14] = 16'hFFFF;  // Neuron 14
    neuron_patterns[ 15] = 16'hFFFF;  // Neuron 15
    neuron_patterns[ 16] = 16'hFFFF;  // Neuron 16
    neuron_patterns[ 17] = 16'hFFFF;  // Neuron 17
    neuron_patterns[ 18] = 16'hFFFF;  // Neuron 18
    neuron_patterns[ 19] = 16'hFFFF;  // Neuron 19
    neuron_patterns[ 20] = 16'hFFFF;  // Neuron 20
    neuron_patterns[ 21] = 16'hFFFF;  // Neuron 21
    neuron_patterns[ 22] = 16'hFFFF;  // Neuron 22
    neuron_patterns[ 23] = 16'hFFFF;  // Neuron 23
    neuron_patterns[ 24] = 16'hFFFF;  // Neuron 24
    neuron_patterns[ 25] = 16'hFFFF;  // Neuron 25
    neuron_patterns[ 26] = 16'hFFFF;  // Neuron 26
    neuron_patterns[ 27] = 16'hFFFF;  // Neuron 27
    neuron_patterns[ 28] = 16'hFFFF;  // Neuron 28
    neuron_patterns[ 29] = 16'hFFFF;  // Neuron 29
    neuron_patterns[ 30] = 16'hFFFF;  // Neuron 30
    neuron_patterns[ 31] = 16'hFFFF;  // Neuron 31
    neuron_patterns[ 32] = 16'hFFFF;  // Neuron 32
    neuron_patterns[ 33] = 16'hFFFF;  // Neuron 33
    neuron_patterns[ 34] = 16'hFFFF;  // Neuron 34
    neuron_patterns[ 35] = 16'hFFFF;  // Neuron 35
    neuron_patterns[ 36] = 16'hFFFF;  // Neuron 36
    neuron_patterns[ 37] = 16'hFFFF;  // Neuron 37
    neuron_patterns[ 38] = 16'hFFFF;  // Neuron 38
    neuron_patterns[ 39] = 16'hFFFF;  // Neuron 39
    neuron_patterns[ 40] = 16'hFFFF;  // Neuron 40
    neuron_patterns[ 41] = 16'hFFFF;  // Neuron 41
    neuron_patterns[ 42] = 16'hFFFF;  // Neuron 42
    neuron_patterns[ 43] = 16'hFFFF;  // Neuron 43
    neuron_patterns[ 44] = 16'hFFFF;  // Neuron 44
    neuron_patterns[ 45] = 16'hFFFF;  // Neuron 45
    neuron_patterns[ 46] = 16'hFFFF;  // Neuron 46
    neuron_patterns[ 47] = 16'hFFFF;  // Neuron 47
    neuron_patterns[ 48] = 16'hFFFF;  // Neuron 48
    neuron_patterns[ 49] = 16'hFFFF;  // Neuron 49
    neuron_patterns[ 50] = 16'hFFFF;  // Neuron 50
    neuron_patterns[ 51] = 16'hFFFF;  // Neuron 51
    neuron_patterns[ 52] = 16'hFFFF;  // Neuron 52
    neuron_patterns[ 53] = 16'hFFFF;  // Neuron 53
    neuron_patterns[ 54] = 16'hFFFF;  // Neuron 54
    neuron_patterns[ 55] = 16'hFFFF;  // Neuron 55
    neuron_patterns[ 56] = 16'hFFFF;  // Neuron 56
    neuron_patterns[ 57] = 16'hFFFF;  // Neuron 57
    neuron_patterns[ 58] = 16'hFFFF;  // Neuron 58
    neuron_patterns[ 59] = 16'hFFFF;  // Neuron 59
    neuron_patterns[ 60] = 16'hFFFF;  // Neuron 60
    neuron_patterns[ 61] = 16'hFFFF;  // Neuron 61
    neuron_patterns[ 62] = 16'hFFFF;  // Neuron 62
    neuron_patterns[ 63] = 16'hFFFF;  // Neuron 63
    neuron_patterns[ 64] = 16'hFFFF;  // Neuron 64
    neuron_patterns[ 65] = 16'hFFFF;  // Neuron 65
    neuron_patterns[ 66] = 16'hFFFF;  // Neuron 66
    neuron_patterns[ 67] = 16'hFFFF;  // Neuron 67
    neuron_patterns[ 68] = 16'hFFFF;  // Neuron 68
    neuron_patterns[ 69] = 16'hFFFF;  // Neuron 69
    neuron_patterns[ 70] = 16'hFFFF;  // Neuron 70
    neuron_patterns[ 71] = 16'hFFFF;  // Neuron 71
    neuron_patterns[ 72] = 16'hFFFF;  // Neuron 72
    neuron_patterns[ 73] = 16'hFFFF;  // Neuron 73
    neuron_patterns[ 74] = 16'hFFFF;  // Neuron 74
    neuron_patterns[ 75] = 16'hFFFF;  // Neuron 75
    neuron_patterns[ 76] = 16'hFFFF;  // Neuron 76
    neuron_patterns[ 77] = 16'hFFFF;  // Neuron 77
    neuron_patterns[ 78] = 16'hFFFF;  // Neuron 78
    neuron_patterns[ 79] = 16'hFFFF;  // Neuron 79
    neuron_patterns[ 80] = 16'hFFFF;  // Neuron 80
    neuron_patterns[ 81] = 16'hFFFF;  // Neuron 81
    neuron_patterns[ 82] = 16'hFFFF;  // Neuron 82
    neuron_patterns[ 83] = 16'hFFFF;  // Neuron 83
    neuron_patterns[ 84] = 16'hFFFF;  // Neuron 84
    neuron_patterns[ 85] = 16'hFFFF;  // Neuron 85
    neuron_patterns[ 86] = 16'hFFFF;  // Neuron 86
    neuron_patterns[ 87] = 16'hFFFF;  // Neuron 87
    neuron_patterns[ 88] = 16'hFFFF;  // Neuron 88
    neuron_patterns[ 89] = 16'hFFFF;  // Neuron 89
    neuron_patterns[ 90] = 16'hFFFF;  // Neuron 90
    neuron_patterns[ 91] = 16'hFFFF;  // Neuron 91
    neuron_patterns[ 92] = 16'hFFFF;  // Neuron 92
    neuron_patterns[ 93] = 16'hFFFF;  // Neuron 93
    neuron_patterns[ 94] = 16'hFFFF;  // Neuron 94
    neuron_patterns[ 95] = 16'hFFFF;  // Neuron 95
    neuron_patterns[ 96] = 16'hFFFF;  // Neuron 96
    neuron_patterns[ 97] = 16'hFFFF;  // Neuron 97
    neuron_patterns[ 98] = 16'hFFFF;  // Neuron 98
    neuron_patterns[ 99] = 16'hFFFF;  // Neuron 99
    neuron_patterns[100] = 16'hFFFF;  // Neuron 100
    neuron_patterns[101] = 16'hFFFF;  // Neuron 101
    neuron_patterns[102] = 16'hFFFF;  // Neuron 102
    neuron_patterns[103] = 16'hFFFF;  // Neuron 103
    neuron_patterns[104] = 16'hFFFF;  // Neuron 104
    neuron_patterns[105] = 16'hFFFF;  // Neuron 105
    neuron_patterns[106] = 16'hFFFF;  // Neuron 106
    neuron_patterns[107] = 16'hFFFF;  // Neuron 107
    neuron_patterns[108] = 16'hFFFF;  // Neuron 108
    neuron_patterns[109] = 16'hFFFF;  // Neuron 109
    neuron_patterns[110] = 16'hFFFF;  // Neuron 110
    neuron_patterns[111] = 16'hFFFF;  // Neuron 111
    neuron_patterns[112] = 16'hFFFF;  // Neuron 112
    neuron_patterns[113] = 16'hFFFF;  // Neuron 113
    neuron_patterns[114] = 16'hFFFF;  // Neuron 114
    neuron_patterns[115] = 16'hFFFF;  // Neuron 115
    neuron_patterns[116] = 16'hFFFF;  // Neuron 116
    neuron_patterns[117] = 16'hFFFF;  // Neuron 117
    neuron_patterns[118] = 16'hFFFF;  // Neuron 118
    neuron_patterns[119] = 16'hFFFF;  // Neuron 119
    neuron_patterns[120] = 16'hFFFF;  // Neuron 120
    neuron_patterns[121] = 16'hFFFF;  // Neuron 121
    neuron_patterns[122] = 16'hFFFF;  // Neuron 122
    neuron_patterns[123] = 16'hFFFF;  // Neuron 123
    neuron_patterns[124] = 16'hFFFF;  // Neuron 124
    neuron_patterns[125] = 16'hFFFF;  // Neuron 125
    neuron_patterns[126] = 16'hFFFF;  // Neuron 126
    neuron_patterns[127] = 16'hFFFF;  // Neuron 127
    neuron_patterns[128] = 16'hFFFF;  // Neuron 128
    neuron_patterns[129] = 16'hFFFF;  // Neuron 129
    neuron_patterns[130] = 16'hFFFF;  // Neuron 130
    neuron_patterns[131] = 16'hFFFF;  // Neuron 131
    neuron_patterns[132] = 16'hFFFF;  // Neuron 132
    neuron_patterns[133] = 16'hFFFF;  // Neuron 133
    neuron_patterns[134] = 16'hFFFF;  // Neuron 134
    neuron_patterns[135] = 16'hFFFF;  // Neuron 135
    neuron_patterns[136] = 16'hFFFF;  // Neuron 136
    neuron_patterns[137] = 16'hFFFF;  // Neuron 137
    neuron_patterns[138] = 16'hFFFF;  // Neuron 138
    neuron_patterns[139] = 16'hFFFF;  // Neuron 139
    neuron_patterns[140] = 16'hFFFF;  // Neuron 140
    neuron_patterns[141] = 16'hFFFF;  // Neuron 141
    neuron_patterns[142] = 16'hFFFF;  // Neuron 142
    neuron_patterns[143] = 16'hFFFF;  // Neuron 143
    neuron_patterns[144] = 16'hFFFF;  // Neuron 144
    neuron_patterns[145] = 16'hFFFF;  // Neuron 145
    neuron_patterns[146] = 16'hFFFF;  // Neuron 146
    neuron_patterns[147] = 16'hFFFF;  // Neuron 147
    neuron_patterns[148] = 16'hFFFF;  // Neuron 148
    neuron_patterns[149] = 16'hFFFF;  // Neuron 149
    neuron_patterns[150] = 16'hFFFF;  // Neuron 150
    neuron_patterns[151] = 16'hFFFF;  // Neuron 151
    neuron_patterns[152] = 16'hFFFF;  // Neuron 152
    neuron_patterns[153] = 16'hFFFF;  // Neuron 153
    neuron_patterns[154] = 16'hFFFF;  // Neuron 154
    neuron_patterns[155] = 16'hFFFF;  // Neuron 155
    neuron_patterns[156] = 16'hFFFF;  // Neuron 156
    neuron_patterns[157] = 16'hFFFF;  // Neuron 157
    neuron_patterns[158] = 16'hFFFF;  // Neuron 158
    neuron_patterns[159] = 16'hFFFF;  // Neuron 159
    neuron_patterns[160] = 16'hFFFF;  // Neuron 160
    neuron_patterns[161] = 16'hFFFF;  // Neuron 161
    neuron_patterns[162] = 16'hFFFF;  // Neuron 162
    neuron_patterns[163] = 16'hFFFF;  // Neuron 163
    neuron_patterns[164] = 16'hFFFF;  // Neuron 164
    neuron_patterns[165] = 16'hFFFF;  // Neuron 165
    neuron_patterns[166] = 16'hFFFF;  // Neuron 166
    neuron_patterns[167] = 16'hFFFF;  // Neuron 167
    neuron_patterns[168] = 16'hFFFF;  // Neuron 168
    neuron_patterns[169] = 16'hFFFF;  // Neuron 169
    neuron_patterns[170] = 16'hFFFF;  // Neuron 170
    neuron_patterns[171] = 16'hFFFF;  // Neuron 171
    neuron_patterns[172] = 16'hFFFF;  // Neuron 172
    neuron_patterns[173] = 16'hFFFF;  // Neuron 173
    neuron_patterns[174] = 16'hFFFF;  // Neuron 174
    neuron_patterns[175] = 16'hFFFF;  // Neuron 175
    neuron_patterns[176] = 16'hFFFF;  // Neuron 176
    neuron_patterns[177] = 16'hFFFF;  // Neuron 177
    neuron_patterns[178] = 16'hFFFF;  // Neuron 178
    neuron_patterns[179] = 16'hFFFF;  // Neuron 179
    neuron_patterns[180] = 16'hFFFF;  // Neuron 180
    neuron_patterns[181] = 16'hFFFF;  // Neuron 181
    neuron_patterns[182] = 16'hFFFF;  // Neuron 182
    neuron_patterns[183] = 16'hFFFF;  // Neuron 183
    neuron_patterns[184] = 16'hFFFF;  // Neuron 184
    neuron_patterns[185] = 16'hFFFF;  // Neuron 185
    neuron_patterns[186] = 16'hFFFF;  // Neuron 186
    neuron_patterns[187] = 16'hFFFF;  // Neuron 187
    neuron_patterns[188] = 16'hFFFF;  // Neuron 188
    neuron_patterns[189] = 16'hFFFF;  // Neuron 189
    neuron_patterns[190] = 16'hFFFF;  // Neuron 190
    neuron_patterns[191] = 16'hFFFF;  // Neuron 191
    neuron_patterns[192] = 16'hFFFF;  // Neuron 192
    neuron_patterns[193] = 16'hFFFF;  // Neuron 193
    neuron_patterns[194] = 16'hFFFF;  // Neuron 194
    neuron_patterns[195] = 16'hFFFF;  // Neuron 195
    neuron_patterns[196] = 16'hFFFF;  // Neuron 196
    neuron_patterns[197] = 16'hFFFF;  // Neuron 197
    neuron_patterns[198] = 16'hFFFF;  // Neuron 198
    neuron_patterns[199] = 16'hFFFF;  // Neuron 199
    neuron_patterns[200] = 16'hFFFF;  // Neuron 200
    neuron_patterns[201] = 16'hFFFF;  // Neuron 201
    neuron_patterns[202] = 16'hFFFF;  // Neuron 202
    neuron_patterns[203] = 16'hFFFF;  // Neuron 203
    neuron_patterns[204] = 16'hFFFF;  // Neuron 204
    neuron_patterns[205] = 16'hFFFF;  // Neuron 205
    neuron_patterns[206] = 16'hFFFF;  // Neuron 206
    neuron_patterns[207] = 16'hFFFF;  // Neuron 207
    neuron_patterns[208] = 16'hFFFF;  // Neuron 208
    neuron_patterns[209] = 16'hFFFF;  // Neuron 209
    neuron_patterns[210] = 16'hFFFF;  // Neuron 210
    neuron_patterns[211] = 16'hFFFF;  // Neuron 211
    neuron_patterns[212] = 16'hFFFF;  // Neuron 212
    neuron_patterns[213] = 16'hFFFF;  // Neuron 213
    neuron_patterns[214] = 16'hFFFF;  // Neuron 214
    neuron_patterns[215] = 16'hFFFF;  // Neuron 215
    neuron_patterns[216] = 16'hFFFF;  // Neuron 216
    neuron_patterns[217] = 16'hFFFF;  // Neuron 217
    neuron_patterns[218] = 16'hFFFF;  // Neuron 218
    neuron_patterns[219] = 16'hFFFF;  // Neuron 219
    neuron_patterns[220] = 16'hFFFF;  // Neuron 220
    neuron_patterns[221] = 16'hFFFF;  // Neuron 221
    neuron_patterns[222] = 16'hFFFF;  // Neuron 222
    neuron_patterns[223] = 16'hFFFF;  // Neuron 223
    neuron_patterns[224] = 16'hFFFF;  // Neuron 224
    neuron_patterns[225] = 16'hFFFF;  // Neuron 225
    neuron_patterns[226] = 16'hFFFF;  // Neuron 226
    neuron_patterns[227] = 16'hFFFF;  // Neuron 227
    neuron_patterns[228] = 16'hFFFF;  // Neuron 228
    neuron_patterns[229] = 16'hFFFF;  // Neuron 229
    neuron_patterns[230] = 16'hFFFF;  // Neuron 230
    neuron_patterns[231] = 16'hFFFF;  // Neuron 231
    neuron_patterns[232] = 16'hFFFF;  // Neuron 232
    neuron_patterns[233] = 16'hFFFF;  // Neuron 233
    neuron_patterns[234] = 16'hFFFF;  // Neuron 234
    neuron_patterns[235] = 16'hFFFF;  // Neuron 235
    neuron_patterns[236] = 16'hFFFF;  // Neuron 236
    neuron_patterns[237] = 16'hFFFF;  // Neuron 237
    neuron_patterns[238] = 16'hFFFF;  // Neuron 238
    neuron_patterns[239] = 16'hFFFF;  // Neuron 239
    neuron_patterns[240] = 16'hFFFF;  // Neuron 240
    neuron_patterns[241] = 16'hFFFF;  // Neuron 241
    neuron_patterns[242] = 16'hFFFF;  // Neuron 242
    neuron_patterns[243] = 16'hFFFF;  // Neuron 243
    neuron_patterns[244] = 16'hFFFF;  // Neuron 244
    neuron_patterns[245] = 16'hFFFF;  // Neuron 245
    neuron_patterns[246] = 16'hFFFF;  // Neuron 246
    neuron_patterns[247] = 16'hFFFF;  // Neuron 247
    neuron_patterns[248] = 16'hFFFF;  // Neuron 248
    neuron_patterns[249] = 16'hFFFF;  // Neuron 249
    neuron_patterns[250] = 16'hFFFF;  // Neuron 250
    neuron_patterns[251] = 16'hFFFF;  // Neuron 251
    neuron_patterns[252] = 16'hFFFF;  // Neuron 252
    neuron_patterns[253] = 16'hFFFF;  // Neuron 253
    neuron_patterns[254] = 16'hFFFF;  // Neuron 254
    neuron_patterns[255] = 16'hFFFF;  // Neuron 255
  end

endmodule
