// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module attention_enc_10_q_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h1000;
    tile_memory[  1] = 16'h0001;
    tile_memory[  2] = 16'h2001;
    tile_memory[  3] = 16'h0002;
    tile_memory[  4] = 16'h0014;
    tile_memory[  5] = 16'h0901;
    tile_memory[  6] = 16'h0001;
    tile_memory[  7] = 16'h4020;
    tile_memory[  8] = 16'h0040;
    tile_memory[  9] = 16'h001A;
    tile_memory[ 10] = 16'h4400;
    tile_memory[ 11] = 16'h0801;
    tile_memory[ 12] = 16'h0800;
    tile_memory[ 13] = 16'h0200;
    tile_memory[ 14] = 16'h2000;
    tile_memory[ 15] = 16'h8000;
    tile_memory[ 16] = 16'h0041;
    tile_memory[ 17] = 16'h0202;
    tile_memory[ 18] = 16'h0480;
    tile_memory[ 19] = 16'h8000;
    tile_memory[ 20] = 16'h0004;
    tile_memory[ 21] = 16'h0500;
    tile_memory[ 22] = 16'h0002;
    tile_memory[ 23] = 16'h0020;
    tile_memory[ 24] = 16'h0008;
    tile_memory[ 25] = 16'h2000;
    tile_memory[ 26] = 16'h1040;
    tile_memory[ 27] = 16'h0404;
    tile_memory[ 28] = 16'h0400;
    tile_memory[ 29] = 16'h4080;
    tile_memory[ 30] = 16'h1000;
    tile_memory[ 31] = 16'h000A;
    tile_memory[ 32] = 16'h2000;
    tile_memory[ 33] = 16'h0080;
    tile_memory[ 34] = 16'h0006;
    tile_memory[ 35] = 16'h4002;
    tile_memory[ 36] = 16'h0044;
    tile_memory[ 37] = 16'h8800;
    tile_memory[ 38] = 16'h8000;
    tile_memory[ 39] = 16'h0800;
    tile_memory[ 40] = 16'h0020;
    tile_memory[ 41] = 16'h0C00;
    tile_memory[ 42] = 16'h8000;
    tile_memory[ 43] = 16'h2001;
    tile_memory[ 44] = 16'h0020;
    tile_memory[ 45] = 16'h0088;
    tile_memory[ 46] = 16'h2200;
    tile_memory[ 47] = 16'h0002;
    tile_memory[ 48] = 16'h1000;
    tile_memory[ 49] = 16'h2000;
    tile_memory[ 50] = 16'h2001;
    tile_memory[ 51] = 16'h0002;
    tile_memory[ 52] = 16'h0014;
    tile_memory[ 53] = 16'h0901;
    tile_memory[ 54] = 16'h0001;
    tile_memory[ 55] = 16'h4020;
    tile_memory[ 56] = 16'h0040;
    tile_memory[ 57] = 16'h001A;
    tile_memory[ 58] = 16'h4400;
    tile_memory[ 59] = 16'h0801;
    tile_memory[ 60] = 16'h0800;
    tile_memory[ 61] = 16'h0200;
    tile_memory[ 62] = 16'h0040;
    tile_memory[ 63] = 16'h8000;
    tile_memory[ 64] = 16'h0041;
    tile_memory[ 65] = 16'h0801;
    tile_memory[ 66] = 16'h2031;
    tile_memory[ 67] = 16'h0102;
    tile_memory[ 68] = 16'h0214;
    tile_memory[ 69] = 16'h0500;
    tile_memory[ 70] = 16'h1011;
    tile_memory[ 71] = 16'h0020;
    tile_memory[ 72] = 16'h0008;
    tile_memory[ 73] = 16'h2000;
    tile_memory[ 74] = 16'h1040;
    tile_memory[ 75] = 16'h0404;
    tile_memory[ 76] = 16'h0400;
    tile_memory[ 77] = 16'h4080;
    tile_memory[ 78] = 16'h2100;
    tile_memory[ 79] = 16'h8008;
    tile_memory[ 80] = 16'h00C1;
    tile_memory[ 81] = 16'h0382;
    tile_memory[ 82] = 16'h0C80;
    tile_memory[ 83] = 16'h8050;
    tile_memory[ 84] = 16'h0844;
    tile_memory[ 85] = 16'h2520;
    tile_memory[ 86] = 16'h0012;
    tile_memory[ 87] = 16'h00A2;
    tile_memory[ 88] = 16'h100A;
    tile_memory[ 89] = 16'h2081;
    tile_memory[ 90] = 16'h1044;
    tile_memory[ 91] = 16'h2484;
    tile_memory[ 92] = 16'h8400;
    tile_memory[ 93] = 16'h4880;
    tile_memory[ 94] = 16'h1044;
    tile_memory[ 95] = 16'h400A;
    tile_memory[ 96] = 16'h1000;
    tile_memory[ 97] = 16'h0180;
    tile_memory[ 98] = 16'h2001;
    tile_memory[ 99] = 16'h0002;
    tile_memory[100] = 16'h0014;
    tile_memory[101] = 16'h0901;
    tile_memory[102] = 16'h0001;
    tile_memory[103] = 16'h4030;
    tile_memory[104] = 16'h0060;
    tile_memory[105] = 16'h001A;
    tile_memory[106] = 16'h4400;
    tile_memory[107] = 16'h0801;
    tile_memory[108] = 16'h0800;
    tile_memory[109] = 16'h0200;
    tile_memory[110] = 16'h2224;
    tile_memory[111] = 16'h8000;
    tile_memory[112] = 16'h0041;
    tile_memory[113] = 16'hA040;
    tile_memory[114] = 16'h2091;
    tile_memory[115] = 16'h0102;
    tile_memory[116] = 16'h0016;
    tile_memory[117] = 16'h0500;
    tile_memory[118] = 16'h0101;
    tile_memory[119] = 16'h0020;
    tile_memory[120] = 16'h0008;
    tile_memory[121] = 16'h2000;
    tile_memory[122] = 16'h1040;
    tile_memory[123] = 16'h0404;
    tile_memory[124] = 16'h0400;
    tile_memory[125] = 16'h4080;
    tile_memory[126] = 16'h0050;
    tile_memory[127] = 16'h9200;
    tile_memory[128] = 16'h0050;
    tile_memory[129] = 16'h0144;
    tile_memory[130] = 16'h0002;
    tile_memory[131] = 16'h08A0;
    tile_memory[132] = 16'h0088;
    tile_memory[133] = 16'h0A00;
    tile_memory[134] = 16'h0B00;
    tile_memory[135] = 16'h0010;
    tile_memory[136] = 16'h2140;
    tile_memory[137] = 16'h8840;
    tile_memory[138] = 16'h2401;
    tile_memory[139] = 16'h0818;
    tile_memory[140] = 16'h0500;
    tile_memory[141] = 16'h1000;
    tile_memory[142] = 16'h0008;
    tile_memory[143] = 16'h9000;
    tile_memory[144] = 16'h1000;
    tile_memory[145] = 16'h0080;
    tile_memory[146] = 16'h2001;
    tile_memory[147] = 16'h0002;
    tile_memory[148] = 16'h0014;
    tile_memory[149] = 16'h0901;
    tile_memory[150] = 16'h0001;
    tile_memory[151] = 16'h4030;
    tile_memory[152] = 16'h0040;
    tile_memory[153] = 16'h001A;
    tile_memory[154] = 16'h4400;
    tile_memory[155] = 16'h0801;
    tile_memory[156] = 16'h0800;
    tile_memory[157] = 16'h0200;
    tile_memory[158] = 16'h8000;
    tile_memory[159] = 16'h8000;
    tile_memory[160] = 16'h0041;
    tile_memory[161] = 16'hC001;
    tile_memory[162] = 16'h0A02;
    tile_memory[163] = 16'h2040;
    tile_memory[164] = 16'h0040;
    tile_memory[165] = 16'h0500;
    tile_memory[166] = 16'h4018;
    tile_memory[167] = 16'h0020;
    tile_memory[168] = 16'h0008;
    tile_memory[169] = 16'h2000;
    tile_memory[170] = 16'h1040;
    tile_memory[171] = 16'h0404;
    tile_memory[172] = 16'h0400;
    tile_memory[173] = 16'h4080;
    tile_memory[174] = 16'h0008;
    tile_memory[175] = 16'h0002;
    tile_memory[176] = 16'h10A0;
    tile_memory[177] = 16'h1200;
    tile_memory[178] = 16'h2000;
    tile_memory[179] = 16'h010A;
    tile_memory[180] = 16'h4400;
    tile_memory[181] = 16'h2410;
    tile_memory[182] = 16'h000A;
    tile_memory[183] = 16'hC200;
    tile_memory[184] = 16'h0120;
    tile_memory[185] = 16'h0800;
    tile_memory[186] = 16'h8050;
    tile_memory[187] = 16'h0800;
    tile_memory[188] = 16'h8004;
    tile_memory[189] = 16'h4080;
    tile_memory[190] = 16'h0440;
    tile_memory[191] = 16'h0100;
    tile_memory[192] = 16'h1000;
    tile_memory[193] = 16'h3040;
    tile_memory[194] = 16'h2001;
    tile_memory[195] = 16'h0002;
    tile_memory[196] = 16'h0014;
    tile_memory[197] = 16'h0901;
    tile_memory[198] = 16'h0001;
    tile_memory[199] = 16'h4030;
    tile_memory[200] = 16'h0060;
    tile_memory[201] = 16'h001A;
    tile_memory[202] = 16'h4420;
    tile_memory[203] = 16'h0801;
    tile_memory[204] = 16'h0800;
    tile_memory[205] = 16'h0200;
    tile_memory[206] = 16'h0001;
    tile_memory[207] = 16'h8000;
    tile_memory[208] = 16'h0041;
    tile_memory[209] = 16'h2020;
    tile_memory[210] = 16'h3400;
    tile_memory[211] = 16'h0088;
    tile_memory[212] = 16'h8010;
    tile_memory[213] = 16'h0500;
    tile_memory[214] = 16'h1006;
    tile_memory[215] = 16'h0020;
    tile_memory[216] = 16'h0008;
    tile_memory[217] = 16'h2000;
    tile_memory[218] = 16'h1040;
    tile_memory[219] = 16'h0404;
    tile_memory[220] = 16'h0400;
    tile_memory[221] = 16'h4080;
    tile_memory[222] = 16'h0008;
    tile_memory[223] = 16'h0A04;
    tile_memory[224] = 16'h0200;
    tile_memory[225] = 16'h0109;
    tile_memory[226] = 16'h4C00;
    tile_memory[227] = 16'h1400;
    tile_memory[228] = 16'h0240;
    tile_memory[229] = 16'h0288;
    tile_memory[230] = 16'h2804;
    tile_memory[231] = 16'h0008;
    tile_memory[232] = 16'h5020;
    tile_memory[233] = 16'hA001;
    tile_memory[234] = 16'h0020;
    tile_memory[235] = 16'h1001;
    tile_memory[236] = 16'h1000;
    tile_memory[237] = 16'h0010;
    tile_memory[238] = 16'h8000;
    tile_memory[239] = 16'h1000;
    tile_memory[240] = 16'h1000;
    tile_memory[241] = 16'h0220;
    tile_memory[242] = 16'h2001;
    tile_memory[243] = 16'h0002;
    tile_memory[244] = 16'h0014;
    tile_memory[245] = 16'h0901;
    tile_memory[246] = 16'h0001;
    tile_memory[247] = 16'h4030;
    tile_memory[248] = 16'h0040;
    tile_memory[249] = 16'h001A;
    tile_memory[250] = 16'h4400;
    tile_memory[251] = 16'h0801;
    tile_memory[252] = 16'h0800;
    tile_memory[253] = 16'h0200;
    tile_memory[254] = 16'h4500;
    tile_memory[255] = 16'h8000;
  end

endmodule
