// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module fc_v_enc_10_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h0004;  // Neuron 0
    neuron_patterns[  1] = 16'h6DEA;  // Neuron 1
    neuron_patterns[  2] = 16'h0270;  // Neuron 2
    neuron_patterns[  3] = 16'hEE78;  // Neuron 3
    neuron_patterns[  4] = 16'h8AF5;  // Neuron 4
    neuron_patterns[  5] = 16'h8202;  // Neuron 5
    neuron_patterns[  6] = 16'h2110;  // Neuron 6
    neuron_patterns[  7] = 16'h5CA2;  // Neuron 7
    neuron_patterns[  8] = 16'h2460;  // Neuron 8
    neuron_patterns[  9] = 16'h8931;  // Neuron 9
    neuron_patterns[ 10] = 16'h305E;  // Neuron 10
    neuron_patterns[ 11] = 16'h4802;  // Neuron 11
    neuron_patterns[ 12] = 16'h0F80;  // Neuron 12
    neuron_patterns[ 13] = 16'hCBA0;  // Neuron 13
    neuron_patterns[ 14] = 16'h2BD2;  // Neuron 14
    neuron_patterns[ 15] = 16'h5104;  // Neuron 15
    neuron_patterns[ 16] = 16'hED56;  // Neuron 16
    neuron_patterns[ 17] = 16'h280D;  // Neuron 17
    neuron_patterns[ 18] = 16'h6C8C;  // Neuron 18
    neuron_patterns[ 19] = 16'hD858;  // Neuron 19
    neuron_patterns[ 20] = 16'h98CB;  // Neuron 20
    neuron_patterns[ 21] = 16'h5190;  // Neuron 21
    neuron_patterns[ 22] = 16'h0002;  // Neuron 22
    neuron_patterns[ 23] = 16'h292A;  // Neuron 23
    neuron_patterns[ 24] = 16'h181F;  // Neuron 24
    neuron_patterns[ 25] = 16'hCC40;  // Neuron 25
    neuron_patterns[ 26] = 16'hF482;  // Neuron 26
    neuron_patterns[ 27] = 16'h4BEB;  // Neuron 27
    neuron_patterns[ 28] = 16'h4C26;  // Neuron 28
    neuron_patterns[ 29] = 16'h0723;  // Neuron 29
    neuron_patterns[ 30] = 16'h0C10;  // Neuron 30
    neuron_patterns[ 31] = 16'h8A0C;  // Neuron 31
    neuron_patterns[ 32] = 16'h02BE;  // Neuron 32
    neuron_patterns[ 33] = 16'hD43B;  // Neuron 33
    neuron_patterns[ 34] = 16'h1124;  // Neuron 34
    neuron_patterns[ 35] = 16'h941C;  // Neuron 35
    neuron_patterns[ 36] = 16'h0880;  // Neuron 36
    neuron_patterns[ 37] = 16'h8C8C;  // Neuron 37
    neuron_patterns[ 38] = 16'hE267;  // Neuron 38
    neuron_patterns[ 39] = 16'h643D;  // Neuron 39
    neuron_patterns[ 40] = 16'h09F2;  // Neuron 40
    neuron_patterns[ 41] = 16'h4150;  // Neuron 41
    neuron_patterns[ 42] = 16'h8809;  // Neuron 42
    neuron_patterns[ 43] = 16'h0403;  // Neuron 43
    neuron_patterns[ 44] = 16'h0008;  // Neuron 44
    neuron_patterns[ 45] = 16'h73C4;  // Neuron 45
    neuron_patterns[ 46] = 16'h2339;  // Neuron 46
    neuron_patterns[ 47] = 16'h0948;  // Neuron 47
    neuron_patterns[ 48] = 16'h008D;  // Neuron 48
    neuron_patterns[ 49] = 16'h6DAA;  // Neuron 49
    neuron_patterns[ 50] = 16'h2222;  // Neuron 50
    neuron_patterns[ 51] = 16'hCA72;  // Neuron 51
    neuron_patterns[ 52] = 16'h87F0;  // Neuron 52
    neuron_patterns[ 53] = 16'hC882;  // Neuron 53
    neuron_patterns[ 54] = 16'hA140;  // Neuron 54
    neuron_patterns[ 55] = 16'h4CB1;  // Neuron 55
    neuron_patterns[ 56] = 16'h2600;  // Neuron 56
    neuron_patterns[ 57] = 16'h102D;  // Neuron 57
    neuron_patterns[ 58] = 16'hF446;  // Neuron 58
    neuron_patterns[ 59] = 16'h5020;  // Neuron 59
    neuron_patterns[ 60] = 16'h8D00;  // Neuron 60
    neuron_patterns[ 61] = 16'hC081;  // Neuron 61
    neuron_patterns[ 62] = 16'hA874;  // Neuron 62
    neuron_patterns[ 63] = 16'h4406;  // Neuron 63
    neuron_patterns[ 64] = 16'hE1D6;  // Neuron 64
    neuron_patterns[ 65] = 16'h6809;  // Neuron 65
    neuron_patterns[ 66] = 16'h7028;  // Neuron 66
    neuron_patterns[ 67] = 16'hB868;  // Neuron 67
    neuron_patterns[ 68] = 16'hA3DB;  // Neuron 68
    neuron_patterns[ 69] = 16'h4897;  // Neuron 69
    neuron_patterns[ 70] = 16'h8580;  // Neuron 70
    neuron_patterns[ 71] = 16'h5D02;  // Neuron 71
    neuron_patterns[ 72] = 16'hA80A;  // Neuron 72
    neuron_patterns[ 73] = 16'h0257;  // Neuron 73
    neuron_patterns[ 74] = 16'hE28A;  // Neuron 74
    neuron_patterns[ 75] = 16'h09A1;  // Neuron 75
    neuron_patterns[ 76] = 16'hCCAC;  // Neuron 76
    neuron_patterns[ 77] = 16'h118B;  // Neuron 77
    neuron_patterns[ 78] = 16'h6810;  // Neuron 78
    neuron_patterns[ 79] = 16'hAE00;  // Neuron 79
    neuron_patterns[ 80] = 16'h26BE;  // Neuron 80
    neuron_patterns[ 81] = 16'h857A;  // Neuron 81
    neuron_patterns[ 82] = 16'h1110;  // Neuron 82
    neuron_patterns[ 83] = 16'h8015;  // Neuron 83
    neuron_patterns[ 84] = 16'h24B0;  // Neuron 84
    neuron_patterns[ 85] = 16'h848D;  // Neuron 85
    neuron_patterns[ 86] = 16'h912F;  // Neuron 86
    neuron_patterns[ 87] = 16'hA43D;  // Neuron 87
    neuron_patterns[ 88] = 16'h3280;  // Neuron 88
    neuron_patterns[ 89] = 16'h2150;  // Neuron 89
    neuron_patterns[ 90] = 16'hC88A;  // Neuron 90
    neuron_patterns[ 91] = 16'h1803;  // Neuron 91
    neuron_patterns[ 92] = 16'h0208;  // Neuron 92
    neuron_patterns[ 93] = 16'h512C;  // Neuron 93
    neuron_patterns[ 94] = 16'h317C;  // Neuron 94
    neuron_patterns[ 95] = 16'h0C40;  // Neuron 95
    neuron_patterns[ 96] = 16'h0084;  // Neuron 96
    neuron_patterns[ 97] = 16'h6422;  // Neuron 97
    neuron_patterns[ 98] = 16'h0265;  // Neuron 98
    neuron_patterns[ 99] = 16'hCC58;  // Neuron 99
    neuron_patterns[100] = 16'h8EE0;  // Neuron 100
    neuron_patterns[101] = 16'h0802;  // Neuron 101
    neuron_patterns[102] = 16'h3340;  // Neuron 102
    neuron_patterns[103] = 16'h4EA2;  // Neuron 103
    neuron_patterns[104] = 16'h0EE8;  // Neuron 104
    neuron_patterns[105] = 16'h00BB;  // Neuron 105
    neuron_patterns[106] = 16'h324E;  // Neuron 106
    neuron_patterns[107] = 16'h4102;  // Neuron 107
    neuron_patterns[108] = 16'h0C01;  // Neuron 108
    neuron_patterns[109] = 16'h4081;  // Neuron 109
    neuron_patterns[110] = 16'hA890;  // Neuron 110
    neuron_patterns[111] = 16'h4000;  // Neuron 111
    neuron_patterns[112] = 16'hF1D4;  // Neuron 112
    neuron_patterns[113] = 16'h2489;  // Neuron 113
    neuron_patterns[114] = 16'h609C;  // Neuron 114
    neuron_patterns[115] = 16'h9808;  // Neuron 115
    neuron_patterns[116] = 16'hC0CB;  // Neuron 116
    neuron_patterns[117] = 16'h0893;  // Neuron 117
    neuron_patterns[118] = 16'h0400;  // Neuron 118
    neuron_patterns[119] = 16'h291B;  // Neuron 119
    neuron_patterns[120] = 16'h080E;  // Neuron 120
    neuron_patterns[121] = 16'h0040;  // Neuron 121
    neuron_patterns[122] = 16'hE0A2;  // Neuron 122
    neuron_patterns[123] = 16'hA92B;  // Neuron 123
    neuron_patterns[124] = 16'hC424;  // Neuron 124
    neuron_patterns[125] = 16'h2123;  // Neuron 125
    neuron_patterns[126] = 16'h0813;  // Neuron 126
    neuron_patterns[127] = 16'h2214;  // Neuron 127
    neuron_patterns[128] = 16'h46B8;  // Neuron 128
    neuron_patterns[129] = 16'hB431;  // Neuron 129
    neuron_patterns[130] = 16'h1580;  // Neuron 130
    neuron_patterns[131] = 16'h0152;  // Neuron 131
    neuron_patterns[132] = 16'h1C92;  // Neuron 132
    neuron_patterns[133] = 16'h0A68;  // Neuron 133
    neuron_patterns[134] = 16'h04AD;  // Neuron 134
    neuron_patterns[135] = 16'hA45F;  // Neuron 135
    neuron_patterns[136] = 16'h305C;  // Neuron 136
    neuron_patterns[137] = 16'h0951;  // Neuron 137
    neuron_patterns[138] = 16'h0888;  // Neuron 138
    neuron_patterns[139] = 16'h2493;  // Neuron 139
    neuron_patterns[140] = 16'h420B;  // Neuron 140
    neuron_patterns[141] = 16'h7702;  // Neuron 141
    neuron_patterns[142] = 16'h2138;  // Neuron 142
    neuron_patterns[143] = 16'hAC48;  // Neuron 143
    neuron_patterns[144] = 16'h0084;  // Neuron 144
    neuron_patterns[145] = 16'h7D2A;  // Neuron 145
    neuron_patterns[146] = 16'h002A;  // Neuron 146
    neuron_patterns[147] = 16'h4C50;  // Neuron 147
    neuron_patterns[148] = 16'h82E0;  // Neuron 148
    neuron_patterns[149] = 16'h6302;  // Neuron 149
    neuron_patterns[150] = 16'h2100;  // Neuron 150
    neuron_patterns[151] = 16'h4CA2;  // Neuron 151
    neuron_patterns[152] = 16'hC4C0;  // Neuron 152
    neuron_patterns[153] = 16'h0139;  // Neuron 153
    neuron_patterns[154] = 16'h704F;  // Neuron 154
    neuron_patterns[155] = 16'h0000;  // Neuron 155
    neuron_patterns[156] = 16'h0408;  // Neuron 156
    neuron_patterns[157] = 16'h4080;  // Neuron 157
    neuron_patterns[158] = 16'h0910;  // Neuron 158
    neuron_patterns[159] = 16'h4000;  // Neuron 159
    neuron_patterns[160] = 16'hF5D4;  // Neuron 160
    neuron_patterns[161] = 16'h6809;  // Neuron 161
    neuron_patterns[162] = 16'h408C;  // Neuron 162
    neuron_patterns[163] = 16'h9900;  // Neuron 163
    neuron_patterns[164] = 16'hA0CA;  // Neuron 164
    neuron_patterns[165] = 16'h0297;  // Neuron 165
    neuron_patterns[166] = 16'h0000;  // Neuron 166
    neuron_patterns[167] = 16'h290B;  // Neuron 167
    neuron_patterns[168] = 16'h080E;  // Neuron 168
    neuron_patterns[169] = 16'h0200;  // Neuron 169
    neuron_patterns[170] = 16'hE088;  // Neuron 170
    neuron_patterns[171] = 16'h4863;  // Neuron 171
    neuron_patterns[172] = 16'h5824;  // Neuron 172
    neuron_patterns[173] = 16'h0302;  // Neuron 173
    neuron_patterns[174] = 16'h0814;  // Neuron 174
    neuron_patterns[175] = 16'h2204;  // Neuron 175
    neuron_patterns[176] = 16'h46B4;  // Neuron 176
    neuron_patterns[177] = 16'h84E0;  // Neuron 177
    neuron_patterns[178] = 16'h1000;  // Neuron 178
    neuron_patterns[179] = 16'hC414;  // Neuron 179
    neuron_patterns[180] = 16'h1C80;  // Neuron 180
    neuron_patterns[181] = 16'h0DC8;  // Neuron 181
    neuron_patterns[182] = 16'h8067;  // Neuron 182
    neuron_patterns[183] = 16'h8E5D;  // Neuron 183
    neuron_patterns[184] = 16'h0290;  // Neuron 184
    neuron_patterns[185] = 16'h414A;  // Neuron 185
    neuron_patterns[186] = 16'h4CC8;  // Neuron 186
    neuron_patterns[187] = 16'h0453;  // Neuron 187
    neuron_patterns[188] = 16'h400B;  // Neuron 188
    neuron_patterns[189] = 16'h6820;  // Neuron 189
    neuron_patterns[190] = 16'h2128;  // Neuron 190
    neuron_patterns[191] = 16'h0948;  // Neuron 191
    neuron_patterns[192] = 16'h0084;  // Neuron 192
    neuron_patterns[193] = 16'h660A;  // Neuron 193
    neuron_patterns[194] = 16'h002A;  // Neuron 194
    neuron_patterns[195] = 16'h4C50;  // Neuron 195
    neuron_patterns[196] = 16'h8EE2;  // Neuron 196
    neuron_patterns[197] = 16'h8002;  // Neuron 197
    neuron_patterns[198] = 16'h3100;  // Neuron 198
    neuron_patterns[199] = 16'h44A2;  // Neuron 199
    neuron_patterns[200] = 16'h4400;  // Neuron 200
    neuron_patterns[201] = 16'h042D;  // Neuron 201
    neuron_patterns[202] = 16'hB24F;  // Neuron 202
    neuron_patterns[203] = 16'h1100;  // Neuron 203
    neuron_patterns[204] = 16'h0C08;  // Neuron 204
    neuron_patterns[205] = 16'hC080;  // Neuron 205
    neuron_patterns[206] = 16'h0812;  // Neuron 206
    neuron_patterns[207] = 16'h4001;  // Neuron 207
    neuron_patterns[208] = 16'hD154;  // Neuron 208
    neuron_patterns[209] = 16'h2089;  // Neuron 209
    neuron_patterns[210] = 16'h488C;  // Neuron 210
    neuron_patterns[211] = 16'h9888;  // Neuron 211
    neuron_patterns[212] = 16'hA0CE;  // Neuron 212
    neuron_patterns[213] = 16'h023A;  // Neuron 213
    neuron_patterns[214] = 16'h8000;  // Neuron 214
    neuron_patterns[215] = 16'h0902;  // Neuron 215
    neuron_patterns[216] = 16'h800E;  // Neuron 216
    neuron_patterns[217] = 16'h0200;  // Neuron 217
    neuron_patterns[218] = 16'hE08A;  // Neuron 218
    neuron_patterns[219] = 16'h6B61;  // Neuron 219
    neuron_patterns[220] = 16'h44A4;  // Neuron 220
    neuron_patterns[221] = 16'h2183;  // Neuron 221
    neuron_patterns[222] = 16'h0815;  // Neuron 222
    neuron_patterns[223] = 16'h0A10;  // Neuron 223
    neuron_patterns[224] = 16'h22A4;  // Neuron 224
    neuron_patterns[225] = 16'hC078;  // Neuron 225
    neuron_patterns[226] = 16'h1180;  // Neuron 226
    neuron_patterns[227] = 16'h8010;  // Neuron 227
    neuron_patterns[228] = 16'h0C00;  // Neuron 228
    neuron_patterns[229] = 16'h0E8A;  // Neuron 229
    neuron_patterns[230] = 16'h8047;  // Neuron 230
    neuron_patterns[231] = 16'h285D;  // Neuron 231
    neuron_patterns[232] = 16'h0210;  // Neuron 232
    neuron_patterns[233] = 16'h1150;  // Neuron 233
    neuron_patterns[234] = 16'hE888;  // Neuron 234
    neuron_patterns[235] = 16'h00D3;  // Neuron 235
    neuron_patterns[236] = 16'h0108;  // Neuron 236
    neuron_patterns[237] = 16'h6100;  // Neuron 237
    neuron_patterns[238] = 16'h6128;  // Neuron 238
    neuron_patterns[239] = 16'h8940;  // Neuron 239
    neuron_patterns[240] = 16'h0084;  // Neuron 240
    neuron_patterns[241] = 16'hE446;  // Neuron 241
    neuron_patterns[242] = 16'h00A2;  // Neuron 242
    neuron_patterns[243] = 16'h4D50;  // Neuron 243
    neuron_patterns[244] = 16'h8260;  // Neuron 244
    neuron_patterns[245] = 16'h2002;  // Neuron 245
    neuron_patterns[246] = 16'h2900;  // Neuron 246
    neuron_patterns[247] = 16'h3EA6;  // Neuron 247
    neuron_patterns[248] = 16'hC401;  // Neuron 248
    neuron_patterns[249] = 16'h00A5;  // Neuron 249
    neuron_patterns[250] = 16'h514F;  // Neuron 250
    neuron_patterns[251] = 16'h0000;  // Neuron 251
    neuron_patterns[252] = 16'h0418;  // Neuron 252
    neuron_patterns[253] = 16'h7080;  // Neuron 253
    neuron_patterns[254] = 16'h0850;  // Neuron 254
    neuron_patterns[255] = 16'h4206;  // Neuron 255
  end

endmodule
