// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module fc_k_enc_3_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h048E;  // Neuron 0
    neuron_patterns[  1] = 16'h0002;  // Neuron 1
    neuron_patterns[  2] = 16'h6020;  // Neuron 2
    neuron_patterns[  3] = 16'h21A0;  // Neuron 3
    neuron_patterns[  4] = 16'h0000;  // Neuron 4
    neuron_patterns[  5] = 16'h02A4;  // Neuron 5
    neuron_patterns[  6] = 16'h50A3;  // Neuron 6
    neuron_patterns[  7] = 16'hC102;  // Neuron 7
    neuron_patterns[  8] = 16'h0819;  // Neuron 8
    neuron_patterns[  9] = 16'hB000;  // Neuron 9
    neuron_patterns[ 10] = 16'h0000;  // Neuron 10
    neuron_patterns[ 11] = 16'h0080;  // Neuron 11
    neuron_patterns[ 12] = 16'h0021;  // Neuron 12
    neuron_patterns[ 13] = 16'h0308;  // Neuron 13
    neuron_patterns[ 14] = 16'h0848;  // Neuron 14
    neuron_patterns[ 15] = 16'h0080;  // Neuron 15
    neuron_patterns[ 16] = 16'hE510;  // Neuron 16
    neuron_patterns[ 17] = 16'h9091;  // Neuron 17
    neuron_patterns[ 18] = 16'h4128;  // Neuron 18
    neuron_patterns[ 19] = 16'h4A03;  // Neuron 19
    neuron_patterns[ 20] = 16'h0402;  // Neuron 20
    neuron_patterns[ 21] = 16'h5000;  // Neuron 21
    neuron_patterns[ 22] = 16'h2883;  // Neuron 22
    neuron_patterns[ 23] = 16'h0500;  // Neuron 23
    neuron_patterns[ 24] = 16'h000A;  // Neuron 24
    neuron_patterns[ 25] = 16'h0006;  // Neuron 25
    neuron_patterns[ 26] = 16'h2240;  // Neuron 26
    neuron_patterns[ 27] = 16'h0100;  // Neuron 27
    neuron_patterns[ 28] = 16'h0100;  // Neuron 28
    neuron_patterns[ 29] = 16'h0A00;  // Neuron 29
    neuron_patterns[ 30] = 16'h4081;  // Neuron 30
    neuron_patterns[ 31] = 16'h5902;  // Neuron 31
    neuron_patterns[ 32] = 16'h0018;  // Neuron 32
    neuron_patterns[ 33] = 16'h1000;  // Neuron 33
    neuron_patterns[ 34] = 16'h1008;  // Neuron 34
    neuron_patterns[ 35] = 16'h4200;  // Neuron 35
    neuron_patterns[ 36] = 16'h0001;  // Neuron 36
    neuron_patterns[ 37] = 16'h4308;  // Neuron 37
    neuron_patterns[ 38] = 16'h0018;  // Neuron 38
    neuron_patterns[ 39] = 16'h0061;  // Neuron 39
    neuron_patterns[ 40] = 16'hA510;  // Neuron 40
    neuron_patterns[ 41] = 16'h1410;  // Neuron 41
    neuron_patterns[ 42] = 16'h4020;  // Neuron 42
    neuron_patterns[ 43] = 16'h4201;  // Neuron 43
    neuron_patterns[ 44] = 16'h15A0;  // Neuron 44
    neuron_patterns[ 45] = 16'hB008;  // Neuron 45
    neuron_patterns[ 46] = 16'h0881;  // Neuron 46
    neuron_patterns[ 47] = 16'h5480;  // Neuron 47
    neuron_patterns[ 48] = 16'h048A;  // Neuron 48
    neuron_patterns[ 49] = 16'h2016;  // Neuron 49
    neuron_patterns[ 50] = 16'h2280;  // Neuron 50
    neuron_patterns[ 51] = 16'h0001;  // Neuron 51
    neuron_patterns[ 52] = 16'h0000;  // Neuron 52
    neuron_patterns[ 53] = 16'h4090;  // Neuron 53
    neuron_patterns[ 54] = 16'hC08A;  // Neuron 54
    neuron_patterns[ 55] = 16'h5142;  // Neuron 55
    neuron_patterns[ 56] = 16'h4009;  // Neuron 56
    neuron_patterns[ 57] = 16'h1021;  // Neuron 57
    neuron_patterns[ 58] = 16'h0080;  // Neuron 58
    neuron_patterns[ 59] = 16'h0200;  // Neuron 59
    neuron_patterns[ 60] = 16'h0000;  // Neuron 60
    neuron_patterns[ 61] = 16'h014C;  // Neuron 61
    neuron_patterns[ 62] = 16'h1050;  // Neuron 62
    neuron_patterns[ 63] = 16'h0020;  // Neuron 63
    neuron_patterns[ 64] = 16'h6510;  // Neuron 64
    neuron_patterns[ 65] = 16'h0410;  // Neuron 65
    neuron_patterns[ 66] = 16'h7528;  // Neuron 66
    neuron_patterns[ 67] = 16'h4204;  // Neuron 67
    neuron_patterns[ 68] = 16'h1420;  // Neuron 68
    neuron_patterns[ 69] = 16'hB000;  // Neuron 69
    neuron_patterns[ 70] = 16'h0080;  // Neuron 70
    neuron_patterns[ 71] = 16'h0481;  // Neuron 71
    neuron_patterns[ 72] = 16'h448A;  // Neuron 72
    neuron_patterns[ 73] = 16'h2016;  // Neuron 73
    neuron_patterns[ 74] = 16'h2384;  // Neuron 74
    neuron_patterns[ 75] = 16'h0863;  // Neuron 75
    neuron_patterns[ 76] = 16'h4A40;  // Neuron 76
    neuron_patterns[ 77] = 16'h1934;  // Neuron 77
    neuron_patterns[ 78] = 16'h408A;  // Neuron 78
    neuron_patterns[ 79] = 16'h51C2;  // Neuron 79
    neuron_patterns[ 80] = 16'h0248;  // Neuron 80
    neuron_patterns[ 81] = 16'h1000;  // Neuron 81
    neuron_patterns[ 82] = 16'h1022;  // Neuron 82
    neuron_patterns[ 83] = 16'h4220;  // Neuron 83
    neuron_patterns[ 84] = 16'h05A1;  // Neuron 84
    neuron_patterns[ 85] = 16'h010C;  // Neuron 85
    neuron_patterns[ 86] = 16'h4024;  // Neuron 86
    neuron_patterns[ 87] = 16'h0080;  // Neuron 87
    neuron_patterns[ 88] = 16'hAD10;  // Neuron 88
    neuron_patterns[ 89] = 16'h8110;  // Neuron 89
    neuron_patterns[ 90] = 16'h5120;  // Neuron 90
    neuron_patterns[ 91] = 16'h4205;  // Neuron 91
    neuron_patterns[ 92] = 16'h14A8;  // Neuron 92
    neuron_patterns[ 93] = 16'h1811;  // Neuron 93
    neuron_patterns[ 94] = 16'h2181;  // Neuron 94
    neuron_patterns[ 95] = 16'h0481;  // Neuron 95
    neuron_patterns[ 96] = 16'h440E;  // Neuron 96
    neuron_patterns[ 97] = 16'h2092;  // Neuron 97
    neuron_patterns[ 98] = 16'h6284;  // Neuron 98
    neuron_patterns[ 99] = 16'h8020;  // Neuron 99
    neuron_patterns[100] = 16'h0100;  // Neuron 100
    neuron_patterns[101] = 16'h4215;  // Neuron 101
    neuron_patterns[102] = 16'h44CB;  // Neuron 102
    neuron_patterns[103] = 16'hC1C2;  // Neuron 103
    neuron_patterns[104] = 16'h4A19;  // Neuron 104
    neuron_patterns[105] = 16'h1042;  // Neuron 105
    neuron_patterns[106] = 16'h4084;  // Neuron 106
    neuron_patterns[107] = 16'h42A2;  // Neuron 107
    neuron_patterns[108] = 16'h80A9;  // Neuron 108
    neuron_patterns[109] = 16'h010C;  // Neuron 109
    neuron_patterns[110] = 16'h01B0;  // Neuron 110
    neuron_patterns[111] = 16'h0011;  // Neuron 111
    neuron_patterns[112] = 16'hE510;  // Neuron 112
    neuron_patterns[113] = 16'h4010;  // Neuron 113
    neuron_patterns[114] = 16'h5124;  // Neuron 114
    neuron_patterns[115] = 16'h4305;  // Neuron 115
    neuron_patterns[116] = 16'h94A0;  // Neuron 116
    neuron_patterns[117] = 16'h9811;  // Neuron 117
    neuron_patterns[118] = 16'hA080;  // Neuron 118
    neuron_patterns[119] = 16'h04C1;  // Neuron 119
    neuron_patterns[120] = 16'h108C;  // Neuron 120
    neuron_patterns[121] = 16'h2EC2;  // Neuron 121
    neuron_patterns[122] = 16'h6214;  // Neuron 122
    neuron_patterns[123] = 16'h00A0;  // Neuron 123
    neuron_patterns[124] = 16'h4850;  // Neuron 124
    neuron_patterns[125] = 16'h0094;  // Neuron 125
    neuron_patterns[126] = 16'h5481;  // Neuron 126
    neuron_patterns[127] = 16'hD0C2;  // Neuron 127
    neuron_patterns[128] = 16'h0218;  // Neuron 128
    neuron_patterns[129] = 16'h3820;  // Neuron 129
    neuron_patterns[130] = 16'h4080;  // Neuron 130
    neuron_patterns[131] = 16'h0A80;  // Neuron 131
    neuron_patterns[132] = 16'h0020;  // Neuron 132
    neuron_patterns[133] = 16'h010C;  // Neuron 133
    neuron_patterns[134] = 16'h0060;  // Neuron 134
    neuron_patterns[135] = 16'h2110;  // Neuron 135
    neuron_patterns[136] = 16'hE510;  // Neuron 136
    neuron_patterns[137] = 16'h0010;  // Neuron 137
    neuron_patterns[138] = 16'h4520;  // Neuron 138
    neuron_patterns[139] = 16'h4605;  // Neuron 139
    neuron_patterns[140] = 16'h1462;  // Neuron 140
    neuron_patterns[141] = 16'h4140;  // Neuron 141
    neuron_patterns[142] = 16'h2080;  // Neuron 142
    neuron_patterns[143] = 16'h0400;  // Neuron 143
    neuron_patterns[144] = 16'h0482;  // Neuron 144
    neuron_patterns[145] = 16'h0462;  // Neuron 145
    neuron_patterns[146] = 16'h3390;  // Neuron 146
    neuron_patterns[147] = 16'h4310;  // Neuron 147
    neuron_patterns[148] = 16'h5010;  // Neuron 148
    neuron_patterns[149] = 16'h0036;  // Neuron 149
    neuron_patterns[150] = 16'h84A1;  // Neuron 150
    neuron_patterns[151] = 16'hD182;  // Neuron 151
    neuron_patterns[152] = 16'h2219;  // Neuron 152
    neuron_patterns[153] = 16'hB040;  // Neuron 153
    neuron_patterns[154] = 16'h4040;  // Neuron 154
    neuron_patterns[155] = 16'h4200;  // Neuron 155
    neuron_patterns[156] = 16'h0080;  // Neuron 156
    neuron_patterns[157] = 16'h0108;  // Neuron 157
    neuron_patterns[158] = 16'h0020;  // Neuron 158
    neuron_patterns[159] = 16'h0300;  // Neuron 159
    neuron_patterns[160] = 16'h65B0;  // Neuron 160
    neuron_patterns[161] = 16'h5010;  // Neuron 161
    neuron_patterns[162] = 16'h4600;  // Neuron 162
    neuron_patterns[163] = 16'h4212;  // Neuron 163
    neuron_patterns[164] = 16'h0400;  // Neuron 164
    neuron_patterns[165] = 16'h1104;  // Neuron 165
    neuron_patterns[166] = 16'h8080;  // Neuron 166
    neuron_patterns[167] = 16'h0001;  // Neuron 167
    neuron_patterns[168] = 16'h4406;  // Neuron 168
    neuron_patterns[169] = 16'h0C22;  // Neuron 169
    neuron_patterns[170] = 16'h71A0;  // Neuron 170
    neuron_patterns[171] = 16'h2181;  // Neuron 171
    neuron_patterns[172] = 16'h1810;  // Neuron 172
    neuron_patterns[173] = 16'h0104;  // Neuron 173
    neuron_patterns[174] = 16'h4081;  // Neuron 174
    neuron_patterns[175] = 16'hC102;  // Neuron 175
    neuron_patterns[176] = 16'h241A;  // Neuron 176
    neuron_patterns[177] = 16'h9800;  // Neuron 177
    neuron_patterns[178] = 16'h0040;  // Neuron 178
    neuron_patterns[179] = 16'h0200;  // Neuron 179
    neuron_patterns[180] = 16'h2009;  // Neuron 180
    neuron_patterns[181] = 16'hC008;  // Neuron 181
    neuron_patterns[182] = 16'h0820;  // Neuron 182
    neuron_patterns[183] = 16'h0530;  // Neuron 183
    neuron_patterns[184] = 16'hE510;  // Neuron 184
    neuron_patterns[185] = 16'h3014;  // Neuron 185
    neuron_patterns[186] = 16'h4328;  // Neuron 186
    neuron_patterns[187] = 16'h4808;  // Neuron 187
    neuron_patterns[188] = 16'h1C20;  // Neuron 188
    neuron_patterns[189] = 16'h5008;  // Neuron 189
    neuron_patterns[190] = 16'hA891;  // Neuron 190
    neuron_patterns[191] = 16'h1444;  // Neuron 191
    neuron_patterns[192] = 16'h1602;  // Neuron 192
    neuron_patterns[193] = 16'h0022;  // Neuron 193
    neuron_patterns[194] = 16'h20A1;  // Neuron 194
    neuron_patterns[195] = 16'h21A1;  // Neuron 195
    neuron_patterns[196] = 16'h0000;  // Neuron 196
    neuron_patterns[197] = 16'h0818;  // Neuron 197
    neuron_patterns[198] = 16'h528B;  // Neuron 198
    neuron_patterns[199] = 16'hD982;  // Neuron 199
    neuron_patterns[200] = 16'h0A1B;  // Neuron 200
    neuron_patterns[201] = 16'h1010;  // Neuron 201
    neuron_patterns[202] = 16'h0000;  // Neuron 202
    neuron_patterns[203] = 16'h0A20;  // Neuron 203
    neuron_patterns[204] = 16'h0021;  // Neuron 204
    neuron_patterns[205] = 16'h0308;  // Neuron 205
    neuron_patterns[206] = 16'h4866;  // Neuron 206
    neuron_patterns[207] = 16'h1000;  // Neuron 207
    neuron_patterns[208] = 16'hA510;  // Neuron 208
    neuron_patterns[209] = 16'h9000;  // Neuron 209
    neuron_patterns[210] = 16'h4128;  // Neuron 210
    neuron_patterns[211] = 16'h4204;  // Neuron 211
    neuron_patterns[212] = 16'h3520;  // Neuron 212
    neuron_patterns[213] = 16'h7009;  // Neuron 213
    neuron_patterns[214] = 16'h0880;  // Neuron 214
    neuron_patterns[215] = 16'h0505;  // Neuron 215
    neuron_patterns[216] = 16'h880A;  // Neuron 216
    neuron_patterns[217] = 16'h2062;  // Neuron 217
    neuron_patterns[218] = 16'h2020;  // Neuron 218
    neuron_patterns[219] = 16'h03A1;  // Neuron 219
    neuron_patterns[220] = 16'h5000;  // Neuron 220
    neuron_patterns[221] = 16'h8810;  // Neuron 221
    neuron_patterns[222] = 16'h50AB;  // Neuron 222
    neuron_patterns[223] = 16'h8942;  // Neuron 223
    neuron_patterns[224] = 16'h0C1D;  // Neuron 224
    neuron_patterns[225] = 16'h1804;  // Neuron 225
    neuron_patterns[226] = 16'h0000;  // Neuron 226
    neuron_patterns[227] = 16'h0200;  // Neuron 227
    neuron_patterns[228] = 16'h0481;  // Neuron 228
    neuron_patterns[229] = 16'hC308;  // Neuron 229
    neuron_patterns[230] = 16'h4826;  // Neuron 230
    neuron_patterns[231] = 16'h0002;  // Neuron 231
    neuron_patterns[232] = 16'hE510;  // Neuron 232
    neuron_patterns[233] = 16'h9710;  // Neuron 233
    neuron_patterns[234] = 16'h4320;  // Neuron 234
    neuron_patterns[235] = 16'h4645;  // Neuron 235
    neuron_patterns[236] = 16'h2520;  // Neuron 236
    neuron_patterns[237] = 16'h7009;  // Neuron 237
    neuron_patterns[238] = 16'h8882;  // Neuron 238
    neuron_patterns[239] = 16'h00E4;  // Neuron 239
    neuron_patterns[240] = 16'h048A;  // Neuron 240
    neuron_patterns[241] = 16'h2222;  // Neuron 241
    neuron_patterns[242] = 16'h22A0;  // Neuron 242
    neuron_patterns[243] = 16'h07A0;  // Neuron 243
    neuron_patterns[244] = 16'h4000;  // Neuron 244
    neuron_patterns[245] = 16'h0081;  // Neuron 245
    neuron_patterns[246] = 16'h0483;  // Neuron 246
    neuron_patterns[247] = 16'hC142;  // Neuron 247
    neuron_patterns[248] = 16'h040C;  // Neuron 248
    neuron_patterns[249] = 16'h1044;  // Neuron 249
    neuron_patterns[250] = 16'h8000;  // Neuron 250
    neuron_patterns[251] = 16'h4202;  // Neuron 251
    neuron_patterns[252] = 16'h0401;  // Neuron 252
    neuron_patterns[253] = 16'h410C;  // Neuron 253
    neuron_patterns[254] = 16'h0864;  // Neuron 254
    neuron_patterns[255] = 16'h0000;  // Neuron 255
  end

endmodule
