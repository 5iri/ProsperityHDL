// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module fc_1_enc_3_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h04E0;  // Neuron 0
    neuron_patterns[  1] = 16'h69F8;  // Neuron 1
    neuron_patterns[  2] = 16'h5EFA;  // Neuron 2
    neuron_patterns[  3] = 16'hE22B;  // Neuron 3
    neuron_patterns[  4] = 16'h8E97;  // Neuron 4
    neuron_patterns[  5] = 16'h86B9;  // Neuron 5
    neuron_patterns[  6] = 16'hC211;  // Neuron 6
    neuron_patterns[  7] = 16'hF0AC;  // Neuron 7
    neuron_patterns[  8] = 16'h3950;  // Neuron 8
    neuron_patterns[  9] = 16'hD931;  // Neuron 9
    neuron_patterns[ 10] = 16'h4077;  // Neuron 10
    neuron_patterns[ 11] = 16'hF92B;  // Neuron 11
    neuron_patterns[ 12] = 16'h3AC2;  // Neuron 12
    neuron_patterns[ 13] = 16'hDB04;  // Neuron 13
    neuron_patterns[ 14] = 16'h6FD2;  // Neuron 14
    neuron_patterns[ 15] = 16'h90E4;  // Neuron 15
    neuron_patterns[ 16] = 16'hFF13;  // Neuron 16
    neuron_patterns[ 17] = 16'h0135;  // Neuron 17
    neuron_patterns[ 18] = 16'hE294;  // Neuron 18
    neuron_patterns[ 19] = 16'h66F3;  // Neuron 19
    neuron_patterns[ 20] = 16'h1A60;  // Neuron 20
    neuron_patterns[ 21] = 16'hF596;  // Neuron 21
    neuron_patterns[ 22] = 16'h0702;  // Neuron 22
    neuron_patterns[ 23] = 16'h3E0D;  // Neuron 23
    neuron_patterns[ 24] = 16'h4851;  // Neuron 24
    neuron_patterns[ 25] = 16'h8941;  // Neuron 25
    neuron_patterns[ 26] = 16'h1C01;  // Neuron 26
    neuron_patterns[ 27] = 16'h09CB;  // Neuron 27
    neuron_patterns[ 28] = 16'h44BB;  // Neuron 28
    neuron_patterns[ 29] = 16'h3EA2;  // Neuron 29
    neuron_patterns[ 30] = 16'h9DC9;  // Neuron 30
    neuron_patterns[ 31] = 16'hA12D;  // Neuron 31
    neuron_patterns[ 32] = 16'h40AA;  // Neuron 32
    neuron_patterns[ 33] = 16'hD4F9;  // Neuron 33
    neuron_patterns[ 34] = 16'h0154;  // Neuron 34
    neuron_patterns[ 35] = 16'hD00F;  // Neuron 35
    neuron_patterns[ 36] = 16'h41E0;  // Neuron 36
    neuron_patterns[ 37] = 16'h870D;  // Neuron 37
    neuron_patterns[ 38] = 16'h6342;  // Neuron 38
    neuron_patterns[ 39] = 16'h61B0;  // Neuron 39
    neuron_patterns[ 40] = 16'h30C3;  // Neuron 40
    neuron_patterns[ 41] = 16'hDA9C;  // Neuron 41
    neuron_patterns[ 42] = 16'hEB93;  // Neuron 42
    neuron_patterns[ 43] = 16'hCC01;  // Neuron 43
    neuron_patterns[ 44] = 16'hD940;  // Neuron 44
    neuron_patterns[ 45] = 16'hBB94;  // Neuron 45
    neuron_patterns[ 46] = 16'hCB77;  // Neuron 46
    neuron_patterns[ 47] = 16'h9EDB;  // Neuron 47
    neuron_patterns[ 48] = 16'h9086;  // Neuron 48
    neuron_patterns[ 49] = 16'h6046;  // Neuron 49
    neuron_patterns[ 50] = 16'h9725;  // Neuron 50
    neuron_patterns[ 51] = 16'h6DB0;  // Neuron 51
    neuron_patterns[ 52] = 16'hE16D;  // Neuron 52
    neuron_patterns[ 53] = 16'h5032;  // Neuron 53
    neuron_patterns[ 54] = 16'hB627;  // Neuron 54
    neuron_patterns[ 55] = 16'h1D46;  // Neuron 55
    neuron_patterns[ 56] = 16'hC684;  // Neuron 56
    neuron_patterns[ 57] = 16'h74EB;  // Neuron 57
    neuron_patterns[ 58] = 16'hE617;  // Neuron 58
    neuron_patterns[ 59] = 16'h7B99;  // Neuron 59
    neuron_patterns[ 60] = 16'hD12F;  // Neuron 60
    neuron_patterns[ 61] = 16'h2832;  // Neuron 61
    neuron_patterns[ 62] = 16'hA66E;  // Neuron 62
    neuron_patterns[ 63] = 16'hB2DD;  // Neuron 63
    neuron_patterns[ 64] = 16'h1C31;  // Neuron 64
    neuron_patterns[ 65] = 16'hA5B8;  // Neuron 65
    neuron_patterns[ 66] = 16'h78AC;  // Neuron 66
    neuron_patterns[ 67] = 16'h1CBC;  // Neuron 67
    neuron_patterns[ 68] = 16'h0280;  // Neuron 68
    neuron_patterns[ 69] = 16'h28A4;  // Neuron 69
    neuron_patterns[ 70] = 16'h540F;  // Neuron 70
    neuron_patterns[ 71] = 16'h91AB;  // Neuron 71
    neuron_patterns[ 72] = 16'hA835;  // Neuron 72
    neuron_patterns[ 73] = 16'hA94E;  // Neuron 73
    neuron_patterns[ 74] = 16'hF002;  // Neuron 74
    neuron_patterns[ 75] = 16'hA0EE;  // Neuron 75
    neuron_patterns[ 76] = 16'hB679;  // Neuron 76
    neuron_patterns[ 77] = 16'h18DA;  // Neuron 77
    neuron_patterns[ 78] = 16'h0B92;  // Neuron 78
    neuron_patterns[ 79] = 16'h1FC8;  // Neuron 79
    neuron_patterns[ 80] = 16'hAFCB;  // Neuron 80
    neuron_patterns[ 81] = 16'hF417;  // Neuron 81
    neuron_patterns[ 82] = 16'h9C5D;  // Neuron 82
    neuron_patterns[ 83] = 16'h5018;  // Neuron 83
    neuron_patterns[ 84] = 16'hEACD;  // Neuron 84
    neuron_patterns[ 85] = 16'h0F4E;  // Neuron 85
    neuron_patterns[ 86] = 16'hC44A;  // Neuron 86
    neuron_patterns[ 87] = 16'h9D9F;  // Neuron 87
    neuron_patterns[ 88] = 16'hFA1D;  // Neuron 88
    neuron_patterns[ 89] = 16'hD65E;  // Neuron 89
    neuron_patterns[ 90] = 16'h08C8;  // Neuron 90
    neuron_patterns[ 91] = 16'hA468;  // Neuron 91
    neuron_patterns[ 92] = 16'h98D9;  // Neuron 92
    neuron_patterns[ 93] = 16'h72C9;  // Neuron 93
    neuron_patterns[ 94] = 16'h9582;  // Neuron 94
    neuron_patterns[ 95] = 16'hE9D3;  // Neuron 95
    neuron_patterns[ 96] = 16'h88D0;  // Neuron 96
    neuron_patterns[ 97] = 16'h0582;  // Neuron 97
    neuron_patterns[ 98] = 16'h3B72;  // Neuron 98
    neuron_patterns[ 99] = 16'hEA9E;  // Neuron 99
    neuron_patterns[100] = 16'h151D;  // Neuron 100
    neuron_patterns[101] = 16'h617E;  // Neuron 101
    neuron_patterns[102] = 16'h0623;  // Neuron 102
    neuron_patterns[103] = 16'h312C;  // Neuron 103
    neuron_patterns[104] = 16'h46AA;  // Neuron 104
    neuron_patterns[105] = 16'hC725;  // Neuron 105
    neuron_patterns[106] = 16'h83B4;  // Neuron 106
    neuron_patterns[107] = 16'h19E2;  // Neuron 107
    neuron_patterns[108] = 16'h7320;  // Neuron 108
    neuron_patterns[109] = 16'h31B4;  // Neuron 109
    neuron_patterns[110] = 16'h9390;  // Neuron 110
    neuron_patterns[111] = 16'h6FDE;  // Neuron 111
    neuron_patterns[112] = 16'h8B74;  // Neuron 112
    neuron_patterns[113] = 16'h7264;  // Neuron 113
    neuron_patterns[114] = 16'h0381;  // Neuron 114
    neuron_patterns[115] = 16'h8625;  // Neuron 115
    neuron_patterns[116] = 16'hDE23;  // Neuron 116
    neuron_patterns[117] = 16'h0F79;  // Neuron 117
    neuron_patterns[118] = 16'h6EB4;  // Neuron 118
    neuron_patterns[119] = 16'h235D;  // Neuron 119
    neuron_patterns[120] = 16'hE1E6;  // Neuron 120
    neuron_patterns[121] = 16'hE8C0;  // Neuron 121
    neuron_patterns[122] = 16'hB415;  // Neuron 122
    neuron_patterns[123] = 16'hA966;  // Neuron 123
    neuron_patterns[124] = 16'h78E4;  // Neuron 124
    neuron_patterns[125] = 16'h764E;  // Neuron 125
    neuron_patterns[126] = 16'hD216;  // Neuron 126
    neuron_patterns[127] = 16'hAF64;  // Neuron 127
    neuron_patterns[128] = 16'h9657;  // Neuron 128
    neuron_patterns[129] = 16'h0B31;  // Neuron 129
    neuron_patterns[130] = 16'hB200;  // Neuron 130
    neuron_patterns[131] = 16'hB08E;  // Neuron 131
    neuron_patterns[132] = 16'h86AE;  // Neuron 132
    neuron_patterns[133] = 16'hAE25;  // Neuron 133
    neuron_patterns[134] = 16'h3196;  // Neuron 134
    neuron_patterns[135] = 16'h1735;  // Neuron 135
    neuron_patterns[136] = 16'h546C;  // Neuron 136
    neuron_patterns[137] = 16'h1C4A;  // Neuron 137
    neuron_patterns[138] = 16'h88E3;  // Neuron 138
    neuron_patterns[139] = 16'h3C73;  // Neuron 139
    neuron_patterns[140] = 16'h406C;  // Neuron 140
    neuron_patterns[141] = 16'h7C57;  // Neuron 141
    neuron_patterns[142] = 16'h8894;  // Neuron 142
    neuron_patterns[143] = 16'h8B19;  // Neuron 143
    neuron_patterns[144] = 16'hC45A;  // Neuron 144
    neuron_patterns[145] = 16'hCACD;  // Neuron 145
    neuron_patterns[146] = 16'hF0EE;  // Neuron 146
    neuron_patterns[147] = 16'hE466;  // Neuron 147
    neuron_patterns[148] = 16'hEA3A;  // Neuron 148
    neuron_patterns[149] = 16'h3EF1;  // Neuron 149
    neuron_patterns[150] = 16'h1565;  // Neuron 150
    neuron_patterns[151] = 16'h74E6;  // Neuron 151
    neuron_patterns[152] = 16'hDA4F;  // Neuron 152
    neuron_patterns[153] = 16'hF58A;  // Neuron 153
    neuron_patterns[154] = 16'hDAF8;  // Neuron 154
    neuron_patterns[155] = 16'h5BF0;  // Neuron 155
    neuron_patterns[156] = 16'h3BE5;  // Neuron 156
    neuron_patterns[157] = 16'h174E;  // Neuron 157
    neuron_patterns[158] = 16'hEC17;  // Neuron 158
    neuron_patterns[159] = 16'h7FF7;  // Neuron 159
    neuron_patterns[160] = 16'h1E42;  // Neuron 160
    neuron_patterns[161] = 16'h17F9;  // Neuron 161
    neuron_patterns[162] = 16'hF4DF;  // Neuron 162
    neuron_patterns[163] = 16'h8ABE;  // Neuron 163
    neuron_patterns[164] = 16'h79FF;  // Neuron 164
    neuron_patterns[165] = 16'hEC79;  // Neuron 165
    neuron_patterns[166] = 16'h3723;  // Neuron 166
    neuron_patterns[167] = 16'hD09B;  // Neuron 167
    neuron_patterns[168] = 16'h84BB;  // Neuron 168
    neuron_patterns[169] = 16'hDD6E;  // Neuron 169
    neuron_patterns[170] = 16'h1DAB;  // Neuron 170
    neuron_patterns[171] = 16'hE4C7;  // Neuron 171
    neuron_patterns[172] = 16'hB46B;  // Neuron 172
    neuron_patterns[173] = 16'h94D4;  // Neuron 173
    neuron_patterns[174] = 16'h98D3;  // Neuron 174
    neuron_patterns[175] = 16'h4811;  // Neuron 175
    neuron_patterns[176] = 16'hA01D;  // Neuron 176
    neuron_patterns[177] = 16'h9A5D;  // Neuron 177
    neuron_patterns[178] = 16'h5AF2;  // Neuron 178
    neuron_patterns[179] = 16'hFF8D;  // Neuron 179
    neuron_patterns[180] = 16'hC3BE;  // Neuron 180
    neuron_patterns[181] = 16'h2CF8;  // Neuron 181
    neuron_patterns[182] = 16'h9167;  // Neuron 182
    neuron_patterns[183] = 16'hFBD8;  // Neuron 183
    neuron_patterns[184] = 16'h6B34;  // Neuron 184
    neuron_patterns[185] = 16'h5DEE;  // Neuron 185
    neuron_patterns[186] = 16'hBE4F;  // Neuron 186
    neuron_patterns[187] = 16'hCD67;  // Neuron 187
    neuron_patterns[188] = 16'h1C49;  // Neuron 188
    neuron_patterns[189] = 16'hD0E8;  // Neuron 189
    neuron_patterns[190] = 16'h6CB3;  // Neuron 190
    neuron_patterns[191] = 16'hFB0F;  // Neuron 191
    neuron_patterns[192] = 16'h9E5F;  // Neuron 192
    neuron_patterns[193] = 16'h77F2;  // Neuron 193
    neuron_patterns[194] = 16'h85FB;  // Neuron 194
    neuron_patterns[195] = 16'hE8D7;  // Neuron 195
    neuron_patterns[196] = 16'h4FDF;  // Neuron 196
    neuron_patterns[197] = 16'h8FBF;  // Neuron 197
    neuron_patterns[198] = 16'hCDED;  // Neuron 198
    neuron_patterns[199] = 16'hCFAB;  // Neuron 199
    neuron_patterns[200] = 16'hB3D7;  // Neuron 200
    neuron_patterns[201] = 16'hD31F;  // Neuron 201
    neuron_patterns[202] = 16'h9A6A;  // Neuron 202
    neuron_patterns[203] = 16'h3CF7;  // Neuron 203
    neuron_patterns[204] = 16'hAE2D;  // Neuron 204
    neuron_patterns[205] = 16'hB5B0;  // Neuron 205
    neuron_patterns[206] = 16'h6914;  // Neuron 206
    neuron_patterns[207] = 16'hCEA8;  // Neuron 207
    neuron_patterns[208] = 16'hE2C2;  // Neuron 208
    neuron_patterns[209] = 16'hBBEF;  // Neuron 209
    neuron_patterns[210] = 16'hFD77;  // Neuron 210
    neuron_patterns[211] = 16'h7365;  // Neuron 211
    neuron_patterns[212] = 16'h577E;  // Neuron 212
    neuron_patterns[213] = 16'hFDB1;  // Neuron 213
    neuron_patterns[214] = 16'hEE73;  // Neuron 214
    neuron_patterns[215] = 16'h4CDF;  // Neuron 215
    neuron_patterns[216] = 16'h7883;  // Neuron 216
    neuron_patterns[217] = 16'hFDFD;  // Neuron 217
    neuron_patterns[218] = 16'hEAC9;  // Neuron 218
    neuron_patterns[219] = 16'h6573;  // Neuron 219
    neuron_patterns[220] = 16'h9EF3;  // Neuron 220
    neuron_patterns[221] = 16'hDB7A;  // Neuron 221
    neuron_patterns[222] = 16'h621E;  // Neuron 222
    neuron_patterns[223] = 16'h843D;  // Neuron 223
    neuron_patterns[224] = 16'h627F;  // Neuron 224
    neuron_patterns[225] = 16'h4DC1;  // Neuron 225
    neuron_patterns[226] = 16'hD0CA;  // Neuron 226
    neuron_patterns[227] = 16'h6C7F;  // Neuron 227
    neuron_patterns[228] = 16'h7BFD;  // Neuron 228
    neuron_patterns[229] = 16'hF4CC;  // Neuron 229
    neuron_patterns[230] = 16'h95DD;  // Neuron 230
    neuron_patterns[231] = 16'h4E70;  // Neuron 231
    neuron_patterns[232] = 16'hCB4C;  // Neuron 232
    neuron_patterns[233] = 16'h6F71;  // Neuron 233
    neuron_patterns[234] = 16'h722E;  // Neuron 234
    neuron_patterns[235] = 16'h502F;  // Neuron 235
    neuron_patterns[236] = 16'h22FC;  // Neuron 236
    neuron_patterns[237] = 16'hBF65;  // Neuron 237
    neuron_patterns[238] = 16'h0917;  // Neuron 238
    neuron_patterns[239] = 16'h863E;  // Neuron 239
    neuron_patterns[240] = 16'hD6D8;  // Neuron 240
    neuron_patterns[241] = 16'h41B5;  // Neuron 241
    neuron_patterns[242] = 16'h751C;  // Neuron 242
    neuron_patterns[243] = 16'h1495;  // Neuron 243
    neuron_patterns[244] = 16'h2F75;  // Neuron 244
    neuron_patterns[245] = 16'hF370;  // Neuron 245
    neuron_patterns[246] = 16'h53E8;  // Neuron 246
    neuron_patterns[247] = 16'h94DF;  // Neuron 247
    neuron_patterns[248] = 16'hD603;  // Neuron 248
    neuron_patterns[249] = 16'hFEE6;  // Neuron 249
    neuron_patterns[250] = 16'h2866;  // Neuron 250
    neuron_patterns[251] = 16'h0F86;  // Neuron 251
    neuron_patterns[252] = 16'h7179;  // Neuron 252
    neuron_patterns[253] = 16'h465A;  // Neuron 253
    neuron_patterns[254] = 16'hF71F;  // Neuron 254
    neuron_patterns[255] = 16'h0CE4;  // Neuron 255
  end

endmodule
