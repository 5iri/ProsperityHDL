// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module conv2d_15_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h0800;  // Neuron 0
    neuron_patterns[  1] = 16'h7E7E;  // Neuron 1
    neuron_patterns[  2] = 16'hFEFE;  // Neuron 2
    neuron_patterns[  3] = 16'h70FC;  // Neuron 3
    neuron_patterns[  4] = 16'h0F00;  // Neuron 4
    neuron_patterns[  5] = 16'hCF4F;  // Neuron 5
    neuron_patterns[  6] = 16'hFEFF;  // Neuron 6
    neuron_patterns[  7] = 16'hF0F0;  // Neuron 7
    neuron_patterns[  8] = 16'h0E00;  // Neuron 8
    neuron_patterns[  9] = 16'h6F7F;  // Neuron 9
    neuron_patterns[ 10] = 16'hFEFF;  // Neuron 10
    neuron_patterns[ 11] = 16'h70FE;  // Neuron 11
    neuron_patterns[ 12] = 16'h7E30;  // Neuron 12
    neuron_patterns[ 13] = 16'hFF7F;  // Neuron 13
    neuron_patterns[ 14] = 16'hFFFF;  // Neuron 14
    neuron_patterns[ 15] = 16'h7EFF;  // Neuron 15
    neuron_patterns[ 16] = 16'h7F7C;  // Neuron 16
    neuron_patterns[ 17] = 16'hFFFF;  // Neuron 17
    neuron_patterns[ 18] = 16'hFEFF;  // Neuron 18
    neuron_patterns[ 19] = 16'hFEFE;  // Neuron 19
    neuron_patterns[ 20] = 16'h6EFF;  // Neuron 20
    neuron_patterns[ 21] = 16'hFFFF;  // Neuron 21
    neuron_patterns[ 22] = 16'hFEFF;  // Neuron 22
    neuron_patterns[ 23] = 16'hE0F2;  // Neuron 23
    neuron_patterns[ 24] = 16'h0000;  // Neuron 24
    neuron_patterns[ 25] = 16'h7F07;  // Neuron 25
    neuron_patterns[ 26] = 16'h7E7E;  // Neuron 26
    neuron_patterns[ 27] = 16'h7C7E;  // Neuron 27
    neuron_patterns[ 28] = 16'h0E00;  // Neuron 28
    neuron_patterns[ 29] = 16'h7F7F;  // Neuron 29
    neuron_patterns[ 30] = 16'hFEFF;  // Neuron 30
    neuron_patterns[ 31] = 16'h70FC;  // Neuron 31
    neuron_patterns[ 32] = 16'h83AF;  // Neuron 32
    neuron_patterns[ 33] = 16'hB282;  // Neuron 33
    neuron_patterns[ 34] = 16'hE7FF;  // Neuron 34
    neuron_patterns[ 35] = 16'hFFFF;  // Neuron 35
    neuron_patterns[ 36] = 16'hFF38;  // Neuron 36
    neuron_patterns[ 37] = 16'hFFFF;  // Neuron 37
    neuron_patterns[ 38] = 16'hFFFF;  // Neuron 38
    neuron_patterns[ 39] = 16'h7EFF;  // Neuron 39
    neuron_patterns[ 40] = 16'h3800;  // Neuron 40
    neuron_patterns[ 41] = 16'h0030;  // Neuron 41
    neuron_patterns[ 42] = 16'h0010;  // Neuron 42
    neuron_patterns[ 43] = 16'h000C;  // Neuron 43
    neuron_patterns[ 44] = 16'hFF7F;  // Neuron 44
    neuron_patterns[ 45] = 16'hFFFF;  // Neuron 45
    neuron_patterns[ 46] = 16'hFFFF;  // Neuron 46
    neuron_patterns[ 47] = 16'h7FFF;  // Neuron 47
    neuron_patterns[ 48] = 16'h1C00;  // Neuron 48
    neuron_patterns[ 49] = 16'hFF1F;  // Neuron 49
    neuron_patterns[ 50] = 16'hFFFF;  // Neuron 50
    neuron_patterns[ 51] = 16'h70FE;  // Neuron 51
    neuron_patterns[ 52] = 16'h3000;  // Neuron 52
    neuron_patterns[ 53] = 16'h0000;  // Neuron 53
    neuron_patterns[ 54] = 16'h1C00;  // Neuron 54
    neuron_patterns[ 55] = 16'h001C;  // Neuron 55
    neuron_patterns[ 56] = 16'h0080;  // Neuron 56
    neuron_patterns[ 57] = 16'h0000;  // Neuron 57
    neuron_patterns[ 58] = 16'h0000;  // Neuron 58
    neuron_patterns[ 59] = 16'h0404;  // Neuron 59
    neuron_patterns[ 60] = 16'h7E00;  // Neuron 60
    neuron_patterns[ 61] = 16'hFE7E;  // Neuron 61
    neuron_patterns[ 62] = 16'hFEFE;  // Neuron 62
    neuron_patterns[ 63] = 16'h7CFE;  // Neuron 63
    neuron_patterns[ 64] = 16'h7C30;  // Neuron 64
    neuron_patterns[ 65] = 16'h7C7C;  // Neuron 65
    neuron_patterns[ 66] = 16'hFCFC;  // Neuron 66
    neuron_patterns[ 67] = 16'h3C7C;  // Neuron 67
    neuron_patterns[ 68] = 16'h0000;  // Neuron 68
    neuron_patterns[ 69] = 16'h40C4;  // Neuron 69
    neuron_patterns[ 70] = 16'h1800;  // Neuron 70
    neuron_patterns[ 71] = 16'h041C;  // Neuron 71
    neuron_patterns[ 72] = 16'h7F7F;  // Neuron 72
    neuron_patterns[ 73] = 16'hFF7F;  // Neuron 73
    neuron_patterns[ 74] = 16'hFFFF;  // Neuron 74
    neuron_patterns[ 75] = 16'h7FFE;  // Neuron 75
    neuron_patterns[ 76] = 16'hAE0C;  // Neuron 76
    neuron_patterns[ 77] = 16'hFFFF;  // Neuron 77
    neuron_patterns[ 78] = 16'hFFFF;  // Neuron 78
    neuron_patterns[ 79] = 16'hF0FE;  // Neuron 79
    neuron_patterns[ 80] = 16'h7C00;  // Neuron 80
    neuron_patterns[ 81] = 16'h7E7E;  // Neuron 81
    neuron_patterns[ 82] = 16'h7E7E;  // Neuron 82
    neuron_patterns[ 83] = 16'h7E7E;  // Neuron 83
    neuron_patterns[ 84] = 16'h78FF;  // Neuron 84
    neuron_patterns[ 85] = 16'h7E7E;  // Neuron 85
    neuron_patterns[ 86] = 16'h7E7E;  // Neuron 86
    neuron_patterns[ 87] = 16'h0C7E;  // Neuron 87
    neuron_patterns[ 88] = 16'h7F00;  // Neuron 88
    neuron_patterns[ 89] = 16'h7F7F;  // Neuron 89
    neuron_patterns[ 90] = 16'hFF7F;  // Neuron 90
    neuron_patterns[ 91] = 16'h707E;  // Neuron 91
    neuron_patterns[ 92] = 16'h1E20;  // Neuron 92
    neuron_patterns[ 93] = 16'h7E7F;  // Neuron 93
    neuron_patterns[ 94] = 16'h7E7E;  // Neuron 94
    neuron_patterns[ 95] = 16'h6070;  // Neuron 95
    neuron_patterns[ 96] = 16'h0000;  // Neuron 96
    neuron_patterns[ 97] = 16'h0454;  // Neuron 97
    neuron_patterns[ 98] = 16'h1402;  // Neuron 98
    neuron_patterns[ 99] = 16'h0C1D;  // Neuron 99
    neuron_patterns[100] = 16'h7E64;  // Neuron 100
    neuron_patterns[101] = 16'hFCFE;  // Neuron 101
    neuron_patterns[102] = 16'hFCFC;  // Neuron 102
    neuron_patterns[103] = 16'h7AFE;  // Neuron 103
    neuron_patterns[104] = 16'h0000;  // Neuron 104
    neuron_patterns[105] = 16'h0000;  // Neuron 105
    neuron_patterns[106] = 16'h5400;  // Neuron 106
    neuron_patterns[107] = 16'h041C;  // Neuron 107
    neuron_patterns[108] = 16'h0000;  // Neuron 108
    neuron_patterns[109] = 16'h1C18;  // Neuron 109
    neuron_patterns[110] = 16'h0000;  // Neuron 110
    neuron_patterns[111] = 16'h0000;  // Neuron 111
    neuron_patterns[112] = 16'h3E00;  // Neuron 112
    neuron_patterns[113] = 16'h7E7E;  // Neuron 113
    neuron_patterns[114] = 16'hFEFE;  // Neuron 114
    neuron_patterns[115] = 16'h70FC;  // Neuron 115
    neuron_patterns[116] = 16'h7EB0;  // Neuron 116
    neuron_patterns[117] = 16'h7F7E;  // Neuron 117
    neuron_patterns[118] = 16'h7E7E;  // Neuron 118
    neuron_patterns[119] = 16'h0C3E;  // Neuron 119
    neuron_patterns[120] = 16'h0001;  // Neuron 120
    neuron_patterns[121] = 16'h0000;  // Neuron 121
    neuron_patterns[122] = 16'h0000;  // Neuron 122
    neuron_patterns[123] = 16'h0105;  // Neuron 123
    neuron_patterns[124] = 16'h0000;  // Neuron 124
    neuron_patterns[125] = 16'h0000;  // Neuron 125
    neuron_patterns[126] = 16'h0040;  // Neuron 126
    neuron_patterns[127] = 16'h0000;  // Neuron 127
    neuron_patterns[128] = 16'hFF7E;  // Neuron 128
    neuron_patterns[129] = 16'hFFFF;  // Neuron 129
    neuron_patterns[130] = 16'hFFFF;  // Neuron 130
    neuron_patterns[131] = 16'h7EFF;  // Neuron 131
    neuron_patterns[132] = 16'hFF7E;  // Neuron 132
    neuron_patterns[133] = 16'hFFFF;  // Neuron 133
    neuron_patterns[134] = 16'hFFFF;  // Neuron 134
    neuron_patterns[135] = 16'hFFFF;  // Neuron 135
    neuron_patterns[136] = 16'hFFFF;  // Neuron 136
    neuron_patterns[137] = 16'h646F;  // Neuron 137
    neuron_patterns[138] = 16'hFCFC;  // Neuron 138
    neuron_patterns[139] = 16'h7CFE;  // Neuron 139
    neuron_patterns[140] = 16'h0000;  // Neuron 140
    neuron_patterns[141] = 16'h4000;  // Neuron 141
    neuron_patterns[142] = 16'h0200;  // Neuron 142
    neuron_patterns[143] = 16'h0000;  // Neuron 143
    neuron_patterns[144] = 16'hFFFE;  // Neuron 144
    neuron_patterns[145] = 16'hFFFF;  // Neuron 145
    neuron_patterns[146] = 16'hFFFF;  // Neuron 146
    neuron_patterns[147] = 16'hFFFF;  // Neuron 147
    neuron_patterns[148] = 16'h7F7E;  // Neuron 148
    neuron_patterns[149] = 16'h7F7F;  // Neuron 149
    neuron_patterns[150] = 16'h7F7D;  // Neuron 150
    neuron_patterns[151] = 16'h007F;  // Neuron 151
    neuron_patterns[152] = 16'hFFFF;  // Neuron 152
    neuron_patterns[153] = 16'hFFFF;  // Neuron 153
    neuron_patterns[154] = 16'hFFFF;  // Neuron 154
    neuron_patterns[155] = 16'hFFFF;  // Neuron 155
    neuron_patterns[156] = 16'h7E3E;  // Neuron 156
    neuron_patterns[157] = 16'hFFFF;  // Neuron 157
    neuron_patterns[158] = 16'hFFFE;  // Neuron 158
    neuron_patterns[159] = 16'hFEFF;  // Neuron 159
    neuron_patterns[160] = 16'h1000;  // Neuron 160
    neuron_patterns[161] = 16'h7F7F;  // Neuron 161
    neuron_patterns[162] = 16'h7F7F;  // Neuron 162
    neuron_patterns[163] = 16'h607E;  // Neuron 163
    neuron_patterns[164] = 16'h7F38;  // Neuron 164
    neuron_patterns[165] = 16'hFFFF;  // Neuron 165
    neuron_patterns[166] = 16'hFFFF;  // Neuron 166
    neuron_patterns[167] = 16'hFEFF;  // Neuron 167
    neuron_patterns[168] = 16'hFE7E;  // Neuron 168
    neuron_patterns[169] = 16'hFEFF;  // Neuron 169
    neuron_patterns[170] = 16'hFEFE;  // Neuron 170
    neuron_patterns[171] = 16'hFFFF;  // Neuron 171
    neuron_patterns[172] = 16'hFFFE;  // Neuron 172
    neuron_patterns[173] = 16'hFFFF;  // Neuron 173
    neuron_patterns[174] = 16'hFFFF;  // Neuron 174
    neuron_patterns[175] = 16'hFFFF;  // Neuron 175
    neuron_patterns[176] = 16'hFFFF;  // Neuron 176
    neuron_patterns[177] = 16'hFFFF;  // Neuron 177
    neuron_patterns[178] = 16'hFEFF;  // Neuron 178
    neuron_patterns[179] = 16'hFCFE;  // Neuron 179
    neuron_patterns[180] = 16'h7F01;  // Neuron 180
    neuron_patterns[181] = 16'hFF7F;  // Neuron 181
    neuron_patterns[182] = 16'hFEFF;  // Neuron 182
    neuron_patterns[183] = 16'h3C7E;  // Neuron 183
    neuron_patterns[184] = 16'hFE84;  // Neuron 184
    neuron_patterns[185] = 16'hFEFF;  // Neuron 185
    neuron_patterns[186] = 16'hFFFE;  // Neuron 186
    neuron_patterns[187] = 16'hFCF8;  // Neuron 187
    neuron_patterns[188] = 16'h0000;  // Neuron 188
    neuron_patterns[189] = 16'h0000;  // Neuron 189
    neuron_patterns[190] = 16'h0000;  // Neuron 190
    neuron_patterns[191] = 16'h0000;  // Neuron 191
    neuron_patterns[192] = 16'h1000;  // Neuron 192
    neuron_patterns[193] = 16'h0414;  // Neuron 193
    neuron_patterns[194] = 16'h3C04;  // Neuron 194
    neuron_patterns[195] = 16'h0C1E;  // Neuron 195
    neuron_patterns[196] = 16'h1800;  // Neuron 196
    neuron_patterns[197] = 16'h0000;  // Neuron 197
    neuron_patterns[198] = 16'h6064;  // Neuron 198
    neuron_patterns[199] = 16'h0000;  // Neuron 199
    neuron_patterns[200] = 16'h0000;  // Neuron 200
    neuron_patterns[201] = 16'h0000;  // Neuron 201
    neuron_patterns[202] = 16'h0000;  // Neuron 202
    neuron_patterns[203] = 16'h0000;  // Neuron 203
    neuron_patterns[204] = 16'hFF7C;  // Neuron 204
    neuron_patterns[205] = 16'hFFFF;  // Neuron 205
    neuron_patterns[206] = 16'hFFFF;  // Neuron 206
    neuron_patterns[207] = 16'hFEFF;  // Neuron 207
    neuron_patterns[208] = 16'hBC00;  // Neuron 208
    neuron_patterns[209] = 16'h7EFE;  // Neuron 209
    neuron_patterns[210] = 16'h7F7E;  // Neuron 210
    neuron_patterns[211] = 16'h687E;  // Neuron 211
    neuron_patterns[212] = 16'hFFFF;  // Neuron 212
    neuron_patterns[213] = 16'hFFFF;  // Neuron 213
    neuron_patterns[214] = 16'hFFFF;  // Neuron 214
    neuron_patterns[215] = 16'hFFFF;  // Neuron 215
    neuron_patterns[216] = 16'hFFFF;  // Neuron 216
    neuron_patterns[217] = 16'hFFFF;  // Neuron 217
    neuron_patterns[218] = 16'hFFFF;  // Neuron 218
    neuron_patterns[219] = 16'hFFFF;  // Neuron 219
    neuron_patterns[220] = 16'hFF7E;  // Neuron 220
    neuron_patterns[221] = 16'hFFFF;  // Neuron 221
    neuron_patterns[222] = 16'hFFFF;  // Neuron 222
    neuron_patterns[223] = 16'h7EFF;  // Neuron 223
    neuron_patterns[224] = 16'hFFFF;  // Neuron 224
    neuron_patterns[225] = 16'hFFFF;  // Neuron 225
    neuron_patterns[226] = 16'hFFFF;  // Neuron 226
    neuron_patterns[227] = 16'hFFFF;  // Neuron 227
    neuron_patterns[228] = 16'h7E00;  // Neuron 228
    neuron_patterns[229] = 16'h7E5E;  // Neuron 229
    neuron_patterns[230] = 16'h7C74;  // Neuron 230
    neuron_patterns[231] = 16'h0074;  // Neuron 231
    neuron_patterns[232] = 16'hFF7E;  // Neuron 232
    neuron_patterns[233] = 16'hFFFF;  // Neuron 233
    neuron_patterns[234] = 16'hFFFF;  // Neuron 234
    neuron_patterns[235] = 16'h70FE;  // Neuron 235
    neuron_patterns[236] = 16'h4CFF;  // Neuron 236
    neuron_patterns[237] = 16'hFE7E;  // Neuron 237
    neuron_patterns[238] = 16'hFCFE;  // Neuron 238
    neuron_patterns[239] = 16'h7CFC;  // Neuron 239
    neuron_patterns[240] = 16'hF080;  // Neuron 240
    neuron_patterns[241] = 16'hFCDC;  // Neuron 241
    neuron_patterns[242] = 16'hFCFC;  // Neuron 242
    neuron_patterns[243] = 16'hFEFC;  // Neuron 243
    neuron_patterns[244] = 16'h7C00;  // Neuron 244
    neuron_patterns[245] = 16'h7F7E;  // Neuron 245
    neuron_patterns[246] = 16'hFF7F;  // Neuron 246
    neuron_patterns[247] = 16'h7EFF;  // Neuron 247
    neuron_patterns[248] = 16'h0100;  // Neuron 248
    neuron_patterns[249] = 16'h0008;  // Neuron 249
    neuron_patterns[250] = 16'h5017;  // Neuron 250
    neuron_patterns[251] = 16'h1C3C;  // Neuron 251
    neuron_patterns[252] = 16'h7F20;  // Neuron 252
    neuron_patterns[253] = 16'hFFFF;  // Neuron 253
    neuron_patterns[254] = 16'hFFFF;  // Neuron 254
    neuron_patterns[255] = 16'h60FE;  // Neuron 255
  end

endmodule
