// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module attention_enc_2_q_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h1824;
    tile_memory[  1] = 16'h2802;
    tile_memory[  2] = 16'h0A00;
    tile_memory[  3] = 16'h8203;
    tile_memory[  4] = 16'h00C1;
    tile_memory[  5] = 16'h3211;
    tile_memory[  6] = 16'hC208;
    tile_memory[  7] = 16'h1080;
    tile_memory[  8] = 16'h0082;
    tile_memory[  9] = 16'h2242;
    tile_memory[ 10] = 16'h44A0;
    tile_memory[ 11] = 16'h0640;
    tile_memory[ 12] = 16'hC354;
    tile_memory[ 13] = 16'h2A04;
    tile_memory[ 14] = 16'hA218;
    tile_memory[ 15] = 16'hD055;
    tile_memory[ 16] = 16'h0C39;
    tile_memory[ 17] = 16'h2004;
    tile_memory[ 18] = 16'h8440;
    tile_memory[ 19] = 16'h124D;
    tile_memory[ 20] = 16'h2351;
    tile_memory[ 21] = 16'h0042;
    tile_memory[ 22] = 16'h0E48;
    tile_memory[ 23] = 16'hD085;
    tile_memory[ 24] = 16'h1824;
    tile_memory[ 25] = 16'h2000;
    tile_memory[ 26] = 16'h0200;
    tile_memory[ 27] = 16'h0003;
    tile_memory[ 28] = 16'h80C1;
    tile_memory[ 29] = 16'h1218;
    tile_memory[ 30] = 16'hC219;
    tile_memory[ 31] = 16'h1084;
    tile_memory[ 32] = 16'h0082;
    tile_memory[ 33] = 16'h2044;
    tile_memory[ 34] = 16'h44A1;
    tile_memory[ 35] = 16'h0400;
    tile_memory[ 36] = 16'hC346;
    tile_memory[ 37] = 16'h0004;
    tile_memory[ 38] = 16'hA258;
    tile_memory[ 39] = 16'hD261;
    tile_memory[ 40] = 16'h0311;
    tile_memory[ 41] = 16'h0004;
    tile_memory[ 42] = 16'h8430;
    tile_memory[ 43] = 16'h1049;
    tile_memory[ 44] = 16'h2311;
    tile_memory[ 45] = 16'h10C2;
    tile_memory[ 46] = 16'h1C59;
    tile_memory[ 47] = 16'hC011;
    tile_memory[ 48] = 16'h0804;
    tile_memory[ 49] = 16'hC000;
    tile_memory[ 50] = 16'h0910;
    tile_memory[ 51] = 16'h020B;
    tile_memory[ 52] = 16'h03E1;
    tile_memory[ 53] = 16'hB619;
    tile_memory[ 54] = 16'h4200;
    tile_memory[ 55] = 16'h0494;
    tile_memory[ 56] = 16'h0196;
    tile_memory[ 57] = 16'hA064;
    tile_memory[ 58] = 16'h44A1;
    tile_memory[ 59] = 16'h0482;
    tile_memory[ 60] = 16'hC345;
    tile_memory[ 61] = 16'h4004;
    tile_memory[ 62] = 16'h2218;
    tile_memory[ 63] = 16'h5229;
    tile_memory[ 64] = 16'h0A21;
    tile_memory[ 65] = 16'h018C;
    tile_memory[ 66] = 16'h8508;
    tile_memory[ 67] = 16'h0060;
    tile_memory[ 68] = 16'h2311;
    tile_memory[ 69] = 16'h3082;
    tile_memory[ 70] = 16'h4E59;
    tile_memory[ 71] = 16'hCC85;
    tile_memory[ 72] = 16'h0944;
    tile_memory[ 73] = 16'h0010;
    tile_memory[ 74] = 16'h0E12;
    tile_memory[ 75] = 16'h0289;
    tile_memory[ 76] = 16'h0861;
    tile_memory[ 77] = 16'hA203;
    tile_memory[ 78] = 16'hC219;
    tile_memory[ 79] = 16'h14A0;
    tile_memory[ 80] = 16'h0094;
    tile_memory[ 81] = 16'hA066;
    tile_memory[ 82] = 16'hC000;
    tile_memory[ 83] = 16'h0412;
    tile_memory[ 84] = 16'hDBD5;
    tile_memory[ 85] = 16'h4040;
    tile_memory[ 86] = 16'hA218;
    tile_memory[ 87] = 16'hD27D;
    tile_memory[ 88] = 16'h3E01;
    tile_memory[ 89] = 16'h9505;
    tile_memory[ 90] = 16'h8519;
    tile_memory[ 91] = 16'h1050;
    tile_memory[ 92] = 16'h2310;
    tile_memory[ 93] = 16'h0286;
    tile_memory[ 94] = 16'h4649;
    tile_memory[ 95] = 16'hC181;
    tile_memory[ 96] = 16'h1804;
    tile_memory[ 97] = 16'h8010;
    tile_memory[ 98] = 16'h8F52;
    tile_memory[ 99] = 16'h931A;
    tile_memory[100] = 16'h0165;
    tile_memory[101] = 16'hBA19;
    tile_memory[102] = 16'h4259;
    tile_memory[103] = 16'h9488;
    tile_memory[104] = 16'h0484;
    tile_memory[105] = 16'hAA66;
    tile_memory[106] = 16'h4022;
    tile_memory[107] = 16'h0CA0;
    tile_memory[108] = 16'hC354;
    tile_memory[109] = 16'h0608;
    tile_memory[110] = 16'hA61C;
    tile_memory[111] = 16'h8E7C;
    tile_memory[112] = 16'h2C21;
    tile_memory[113] = 16'h0501;
    tile_memory[114] = 16'h8599;
    tile_memory[115] = 16'h5250;
    tile_memory[116] = 16'h0251;
    tile_memory[117] = 16'h0086;
    tile_memory[118] = 16'h0449;
    tile_memory[119] = 16'hC385;
    tile_memory[120] = 16'h1884;
    tile_memory[121] = 16'h8000;
    tile_memory[122] = 16'h0F10;
    tile_memory[123] = 16'h0703;
    tile_memory[124] = 16'h81C1;
    tile_memory[125] = 16'hB219;
    tile_memory[126] = 16'hC200;
    tile_memory[127] = 16'hD498;
    tile_memory[128] = 16'h2084;
    tile_memory[129] = 16'hA266;
    tile_memory[130] = 16'h4880;
    tile_memory[131] = 16'h0478;
    tile_memory[132] = 16'hC345;
    tile_memory[133] = 16'h0004;
    tile_memory[134] = 16'hA618;
    tile_memory[135] = 16'h5A55;
    tile_memory[136] = 16'h0C09;
    tile_memory[137] = 16'h0404;
    tile_memory[138] = 16'h8581;
    tile_memory[139] = 16'h4241;
    tile_memory[140] = 16'h2351;
    tile_memory[141] = 16'h4002;
    tile_memory[142] = 16'h0C0A;
    tile_memory[143] = 16'hC185;
    tile_memory[144] = 16'h0800;
    tile_memory[145] = 16'h0002;
    tile_memory[146] = 16'h0A52;
    tile_memory[147] = 16'h0A0B;
    tile_memory[148] = 16'h0841;
    tile_memory[149] = 16'hD609;
    tile_memory[150] = 16'h4014;
    tile_memory[151] = 16'h5040;
    tile_memory[152] = 16'h0080;
    tile_memory[153] = 16'h204A;
    tile_memory[154] = 16'hC020;
    tile_memory[155] = 16'h0410;
    tile_memory[156] = 16'h9105;
    tile_memory[157] = 16'h2000;
    tile_memory[158] = 16'h2018;
    tile_memory[159] = 16'h0C50;
    tile_memory[160] = 16'h0011;
    tile_memory[161] = 16'h0014;
    tile_memory[162] = 16'h8100;
    tile_memory[163] = 16'h1001;
    tile_memory[164] = 16'h2060;
    tile_memory[165] = 16'h2082;
    tile_memory[166] = 16'h4018;
    tile_memory[167] = 16'h0001;
    tile_memory[168] = 16'h1204;
    tile_memory[169] = 16'h0002;
    tile_memory[170] = 16'h0A10;
    tile_memory[171] = 16'h0608;
    tile_memory[172] = 16'h4041;
    tile_memory[173] = 16'h2610;
    tile_memory[174] = 16'h0023;
    tile_memory[175] = 16'h1281;
    tile_memory[176] = 16'h0080;
    tile_memory[177] = 16'h2042;
    tile_memory[178] = 16'hC0A0;
    tile_memory[179] = 16'h0CF2;
    tile_memory[180] = 16'hC314;
    tile_memory[181] = 16'h1000;
    tile_memory[182] = 16'hA604;
    tile_memory[183] = 16'h1054;
    tile_memory[184] = 16'h0C19;
    tile_memory[185] = 16'h0004;
    tile_memory[186] = 16'h80C0;
    tile_memory[187] = 16'h1045;
    tile_memory[188] = 16'h2008;
    tile_memory[189] = 16'h2002;
    tile_memory[190] = 16'h0848;
    tile_memory[191] = 16'hC009;
    tile_memory[192] = 16'h1804;
    tile_memory[193] = 16'h2002;
    tile_memory[194] = 16'h0E40;
    tile_memory[195] = 16'h861B;
    tile_memory[196] = 16'h2141;
    tile_memory[197] = 16'h2611;
    tile_memory[198] = 16'h4401;
    tile_memory[199] = 16'h5089;
    tile_memory[200] = 16'h0004;
    tile_memory[201] = 16'h2242;
    tile_memory[202] = 16'hCB20;
    tile_memory[203] = 16'h06F0;
    tile_memory[204] = 16'hC354;
    tile_memory[205] = 16'h1A00;
    tile_memory[206] = 16'hAE18;
    tile_memory[207] = 16'hD255;
    tile_memory[208] = 16'h3C19;
    tile_memory[209] = 16'h2404;
    tile_memory[210] = 16'h81C0;
    tile_memory[211] = 16'h1249;
    tile_memory[212] = 16'h223A;
    tile_memory[213] = 16'h6886;
    tile_memory[214] = 16'h4C48;
    tile_memory[215] = 16'hC501;
    tile_memory[216] = 16'h1A04;
    tile_memory[217] = 16'h0002;
    tile_memory[218] = 16'h0E50;
    tile_memory[219] = 16'h0400;
    tile_memory[220] = 16'h0141;
    tile_memory[221] = 16'h3600;
    tile_memory[222] = 16'h4001;
    tile_memory[223] = 16'h1088;
    tile_memory[224] = 16'h0180;
    tile_memory[225] = 16'h2042;
    tile_memory[226] = 16'h4420;
    tile_memory[227] = 16'h0CF2;
    tile_memory[228] = 16'hC354;
    tile_memory[229] = 16'h2000;
    tile_memory[230] = 16'hA618;
    tile_memory[231] = 16'h5244;
    tile_memory[232] = 16'h0C19;
    tile_memory[233] = 16'h0004;
    tile_memory[234] = 16'h8580;
    tile_memory[235] = 16'h0240;
    tile_memory[236] = 16'h0210;
    tile_memory[237] = 16'h0082;
    tile_memory[238] = 16'h1008;
    tile_memory[239] = 16'hE481;
    tile_memory[240] = 16'h1800;
    tile_memory[241] = 16'h0002;
    tile_memory[242] = 16'h0850;
    tile_memory[243] = 16'h0009;
    tile_memory[244] = 16'h0141;
    tile_memory[245] = 16'hB409;
    tile_memory[246] = 16'h4200;
    tile_memory[247] = 16'h1088;
    tile_memory[248] = 16'h2180;
    tile_memory[249] = 16'hA846;
    tile_memory[250] = 16'hC120;
    tile_memory[251] = 16'h0EF0;
    tile_memory[252] = 16'hC310;
    tile_memory[253] = 16'h0202;
    tile_memory[254] = 16'hA64C;
    tile_memory[255] = 16'h160C;
  end

endmodule
