// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_o_enc_1_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'hF5D1;
    tile_memory[  1] = 16'hF585;
    tile_memory[  2] = 16'h008E;
    tile_memory[  3] = 16'hB46F;
    tile_memory[  4] = 16'h2000;
    tile_memory[  5] = 16'h5400;
    tile_memory[  6] = 16'hBD9B;
    tile_memory[  7] = 16'hE05D;
    tile_memory[  8] = 16'hD7DA;
    tile_memory[  9] = 16'h3987;
    tile_memory[ 10] = 16'h8BBD;
    tile_memory[ 11] = 16'h4BD8;
    tile_memory[ 12] = 16'h8B3E;
    tile_memory[ 13] = 16'h0244;
    tile_memory[ 14] = 16'h8AFF;
    tile_memory[ 15] = 16'h09F6;
    tile_memory[ 16] = 16'h480D;
    tile_memory[ 17] = 16'h0002;
    tile_memory[ 18] = 16'h1A4E;
    tile_memory[ 19] = 16'hA308;
    tile_memory[ 20] = 16'h14C2;
    tile_memory[ 21] = 16'hE488;
    tile_memory[ 22] = 16'hBF5A;
    tile_memory[ 23] = 16'h3E0A;
    tile_memory[ 24] = 16'h6591;
    tile_memory[ 25] = 16'hD585;
    tile_memory[ 26] = 16'h008C;
    tile_memory[ 27] = 16'hB46F;
    tile_memory[ 28] = 16'h2222;
    tile_memory[ 29] = 16'h5C45;
    tile_memory[ 30] = 16'h8D19;
    tile_memory[ 31] = 16'hE00D;
    tile_memory[ 32] = 16'h935A;
    tile_memory[ 33] = 16'h3885;
    tile_memory[ 34] = 16'h8BBD;
    tile_memory[ 35] = 16'h4BD8;
    tile_memory[ 36] = 16'h8B2A;
    tile_memory[ 37] = 16'h0204;
    tile_memory[ 38] = 16'h9AFF;
    tile_memory[ 39] = 16'h19FE;
    tile_memory[ 40] = 16'h480D;
    tile_memory[ 41] = 16'h0002;
    tile_memory[ 42] = 16'h1A6E;
    tile_memory[ 43] = 16'hAB0A;
    tile_memory[ 44] = 16'h16CA;
    tile_memory[ 45] = 16'hE4B8;
    tile_memory[ 46] = 16'h3F4A;
    tile_memory[ 47] = 16'h0C0A;
    tile_memory[ 48] = 16'hE5D1;
    tile_memory[ 49] = 16'hD585;
    tile_memory[ 50] = 16'h008E;
    tile_memory[ 51] = 16'hB40F;
    tile_memory[ 52] = 16'h2222;
    tile_memory[ 53] = 16'h5C45;
    tile_memory[ 54] = 16'h9D99;
    tile_memory[ 55] = 16'hE00D;
    tile_memory[ 56] = 16'h8342;
    tile_memory[ 57] = 16'h3885;
    tile_memory[ 58] = 16'h8BBD;
    tile_memory[ 59] = 16'h4BD8;
    tile_memory[ 60] = 16'h9B3E;
    tile_memory[ 61] = 16'h0244;
    tile_memory[ 62] = 16'h8AFF;
    tile_memory[ 63] = 16'h09FE;
    tile_memory[ 64] = 16'h580D;
    tile_memory[ 65] = 16'h0002;
    tile_memory[ 66] = 16'h1A6E;
    tile_memory[ 67] = 16'hAB0A;
    tile_memory[ 68] = 16'h37C2;
    tile_memory[ 69] = 16'hC4F8;
    tile_memory[ 70] = 16'hBF48;
    tile_memory[ 71] = 16'h0C0A;
    tile_memory[ 72] = 16'h4590;
    tile_memory[ 73] = 16'h8505;
    tile_memory[ 74] = 16'h20CE;
    tile_memory[ 75] = 16'hB66F;
    tile_memory[ 76] = 16'h2000;
    tile_memory[ 77] = 16'h5405;
    tile_memory[ 78] = 16'hFD9B;
    tile_memory[ 79] = 16'hEA5D;
    tile_memory[ 80] = 16'hC142;
    tile_memory[ 81] = 16'h2805;
    tile_memory[ 82] = 16'h8BBD;
    tile_memory[ 83] = 16'h6BD8;
    tile_memory[ 84] = 16'h9B3E;
    tile_memory[ 85] = 16'h0244;
    tile_memory[ 86] = 16'h9AFF;
    tile_memory[ 87] = 16'hD9FE;
    tile_memory[ 88] = 16'h584F;
    tile_memory[ 89] = 16'h0A02;
    tile_memory[ 90] = 16'h1A4E;
    tile_memory[ 91] = 16'hAB08;
    tile_memory[ 92] = 16'h14C2;
    tile_memory[ 93] = 16'hC488;
    tile_memory[ 94] = 16'h3F4A;
    tile_memory[ 95] = 16'h3C0A;
    tile_memory[ 96] = 16'h0190;
    tile_memory[ 97] = 16'h8505;
    tile_memory[ 98] = 16'h208E;
    tile_memory[ 99] = 16'hBC6F;
    tile_memory[100] = 16'h2202;
    tile_memory[101] = 16'h5445;
    tile_memory[102] = 16'hFD1B;
    tile_memory[103] = 16'hEA5D;
    tile_memory[104] = 16'hC742;
    tile_memory[105] = 16'h3887;
    tile_memory[106] = 16'h8BBD;
    tile_memory[107] = 16'h6BD8;
    tile_memory[108] = 16'h9B3E;
    tile_memory[109] = 16'h0244;
    tile_memory[110] = 16'h8AFF;
    tile_memory[111] = 16'h09FE;
    tile_memory[112] = 16'h584F;
    tile_memory[113] = 16'h0E42;
    tile_memory[114] = 16'h124A;
    tile_memory[115] = 16'h2308;
    tile_memory[116] = 16'h14C2;
    tile_memory[117] = 16'hC488;
    tile_memory[118] = 16'hBF4A;
    tile_memory[119] = 16'h0C0A;
    tile_memory[120] = 16'h05D0;
    tile_memory[121] = 16'h8505;
    tile_memory[122] = 16'h008A;
    tile_memory[123] = 16'hB42F;
    tile_memory[124] = 16'h2000;
    tile_memory[125] = 16'h5400;
    tile_memory[126] = 16'hBD19;
    tile_memory[127] = 16'hE01D;
    tile_memory[128] = 16'h8342;
    tile_memory[129] = 16'h2805;
    tile_memory[130] = 16'h8B3D;
    tile_memory[131] = 16'h4BD8;
    tile_memory[132] = 16'h8B28;
    tile_memory[133] = 16'h0244;
    tile_memory[134] = 16'h8AFF;
    tile_memory[135] = 16'h09FE;
    tile_memory[136] = 16'h4808;
    tile_memory[137] = 16'h0002;
    tile_memory[138] = 16'h1A4A;
    tile_memory[139] = 16'h230A;
    tile_memory[140] = 16'h37EA;
    tile_memory[141] = 16'hE498;
    tile_memory[142] = 16'h8D00;
    tile_memory[143] = 16'h0802;
    tile_memory[144] = 16'h45D0;
    tile_memory[145] = 16'h9505;
    tile_memory[146] = 16'h0088;
    tile_memory[147] = 16'hB40A;
    tile_memory[148] = 16'h2000;
    tile_memory[149] = 16'h1400;
    tile_memory[150] = 16'h0023;
    tile_memory[151] = 16'h4008;
    tile_memory[152] = 16'hC342;
    tile_memory[153] = 16'h2805;
    tile_memory[154] = 16'h8BBD;
    tile_memory[155] = 16'h4BD8;
    tile_memory[156] = 16'h8B28;
    tile_memory[157] = 16'h0204;
    tile_memory[158] = 16'h8AFF;
    tile_memory[159] = 16'h19F6;
    tile_memory[160] = 16'h480F;
    tile_memory[161] = 16'h0A02;
    tile_memory[162] = 16'h0A4A;
    tile_memory[163] = 16'h2308;
    tile_memory[164] = 16'h14C2;
    tile_memory[165] = 16'hE488;
    tile_memory[166] = 16'h2D48;
    tile_memory[167] = 16'h0C02;
    tile_memory[168] = 16'h65D0;
    tile_memory[169] = 16'hD505;
    tile_memory[170] = 16'h0088;
    tile_memory[171] = 16'hB40A;
    tile_memory[172] = 16'h2000;
    tile_memory[173] = 16'h5405;
    tile_memory[174] = 16'hBD9B;
    tile_memory[175] = 16'hE05D;
    tile_memory[176] = 16'hD7DA;
    tile_memory[177] = 16'h3987;
    tile_memory[178] = 16'h8BBD;
    tile_memory[179] = 16'h4BD8;
    tile_memory[180] = 16'h8B2E;
    tile_memory[181] = 16'h0244;
    tile_memory[182] = 16'h8AFF;
    tile_memory[183] = 16'h59FE;
    tile_memory[184] = 16'h2000;
    tile_memory[185] = 16'h0002;
    tile_memory[186] = 16'h020E;
    tile_memory[187] = 16'hA348;
    tile_memory[188] = 16'h15C2;
    tile_memory[189] = 16'hE4F8;
    tile_memory[190] = 16'hBF5A;
    tile_memory[191] = 16'h3E0A;
    tile_memory[192] = 16'h45D0;
    tile_memory[193] = 16'hC505;
    tile_memory[194] = 16'h008E;
    tile_memory[195] = 16'hB46F;
    tile_memory[196] = 16'h2222;
    tile_memory[197] = 16'h5C45;
    tile_memory[198] = 16'hBD9B;
    tile_memory[199] = 16'hE05D;
    tile_memory[200] = 16'hD7DA;
    tile_memory[201] = 16'hB987;
    tile_memory[202] = 16'h8BBD;
    tile_memory[203] = 16'hEBD8;
    tile_memory[204] = 16'h8B3E;
    tile_memory[205] = 16'h0244;
    tile_memory[206] = 16'h9AFF;
    tile_memory[207] = 16'h19FE;
    tile_memory[208] = 16'h584F;
    tile_memory[209] = 16'h0802;
    tile_memory[210] = 16'h1A4E;
    tile_memory[211] = 16'hAB08;
    tile_memory[212] = 16'h14EA;
    tile_memory[213] = 16'hC488;
    tile_memory[214] = 16'hBF5A;
    tile_memory[215] = 16'h3C0A;
    tile_memory[216] = 16'h45D0;
    tile_memory[217] = 16'h9505;
    tile_memory[218] = 16'h0088;
    tile_memory[219] = 16'hB40F;
    tile_memory[220] = 16'h2000;
    tile_memory[221] = 16'h5C01;
    tile_memory[222] = 16'hBD9B;
    tile_memory[223] = 16'hE05D;
    tile_memory[224] = 16'hC75A;
    tile_memory[225] = 16'h3887;
    tile_memory[226] = 16'h8BBD;
    tile_memory[227] = 16'h6BD8;
    tile_memory[228] = 16'h8B2E;
    tile_memory[229] = 16'h0244;
    tile_memory[230] = 16'h8A7F;
    tile_memory[231] = 16'h0976;
    tile_memory[232] = 16'h0202;
    tile_memory[233] = 16'h8000;
    tile_memory[234] = 16'h124A;
    tile_memory[235] = 16'h2308;
    tile_memory[236] = 16'h14CA;
    tile_memory[237] = 16'hC488;
    tile_memory[238] = 16'hBF5A;
    tile_memory[239] = 16'h3E0A;
    tile_memory[240] = 16'h65D1;
    tile_memory[241] = 16'hD505;
    tile_memory[242] = 16'h008A;
    tile_memory[243] = 16'hB42F;
    tile_memory[244] = 16'h0020;
    tile_memory[245] = 16'h5401;
    tile_memory[246] = 16'hBD19;
    tile_memory[247] = 16'hE05D;
    tile_memory[248] = 16'h8342;
    tile_memory[249] = 16'h3885;
    tile_memory[250] = 16'h8BBD;
    tile_memory[251] = 16'h6BD8;
    tile_memory[252] = 16'h8B3E;
    tile_memory[253] = 16'h0244;
    tile_memory[254] = 16'h0A75;
    tile_memory[255] = 16'h0946;
  end

endmodule
