// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module attention_enc_1_kv_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h0505;
    tile_memory[  1] = 16'h6624;
    tile_memory[  2] = 16'h4363;
    tile_memory[  3] = 16'hA421;
    tile_memory[  4] = 16'hCCE4;
    tile_memory[  5] = 16'h7FCF;
    tile_memory[  6] = 16'h3677;
    tile_memory[  7] = 16'h482C;
    tile_memory[  8] = 16'hD0D8;
    tile_memory[  9] = 16'h1A9A;
    tile_memory[ 10] = 16'h131B;
    tile_memory[ 11] = 16'h7515;
    tile_memory[ 12] = 16'hEAE7;
    tile_memory[ 13] = 16'h0F8F;
    tile_memory[ 14] = 16'hA7A7;
    tile_memory[ 15] = 16'h5FBD;
    tile_memory[ 16] = 16'hDB5B;
    tile_memory[ 17] = 16'h889A;
    tile_memory[ 18] = 16'h7070;
    tile_memory[ 19] = 16'h0270;
    tile_memory[ 20] = 16'hFA2A;
    tile_memory[ 21] = 16'hF0F8;
    tile_memory[ 22] = 16'h5A3A;
    tile_memory[ 23] = 16'hD3DA;
    tile_memory[ 24] = 16'hCFDD;
    tile_memory[ 25] = 16'h92DF;
    tile_memory[ 26] = 16'h4F93;
    tile_memory[ 27] = 16'h5F5F;
    tile_memory[ 28] = 16'h5353;
    tile_memory[ 29] = 16'hD5D3;
    tile_memory[ 30] = 16'hF5F5;
    tile_memory[ 31] = 16'h01B5;
    tile_memory[ 32] = 16'h8585;
    tile_memory[ 33] = 16'h6724;
    tile_memory[ 34] = 16'h4363;
    tile_memory[ 35] = 16'hF571;
    tile_memory[ 36] = 16'hCDF5;
    tile_memory[ 37] = 16'h7FCF;
    tile_memory[ 38] = 16'h3677;
    tile_memory[ 39] = 16'hC8A8;
    tile_memory[ 40] = 16'hD1D8;
    tile_memory[ 41] = 16'hDBDB;
    tile_memory[ 42] = 16'h93DB;
    tile_memory[ 43] = 16'hF595;
    tile_memory[ 44] = 16'hEAE7;
    tile_memory[ 45] = 16'h2FAF;
    tile_memory[ 46] = 16'hA6A7;
    tile_memory[ 47] = 16'h7DBC;
    tile_memory[ 48] = 16'hDB7B;
    tile_memory[ 49] = 16'h8C9A;
    tile_memory[ 50] = 16'h7C7C;
    tile_memory[ 51] = 16'h0378;
    tile_memory[ 52] = 16'hBB2B;
    tile_memory[ 53] = 16'hB0B8;
    tile_memory[ 54] = 16'hDB9B;
    tile_memory[ 55] = 16'hF3DB;
    tile_memory[ 56] = 16'hEFFD;
    tile_memory[ 57] = 16'hF2FF;
    tile_memory[ 58] = 16'h4FB3;
    tile_memory[ 59] = 16'h5D5D;
    tile_memory[ 60] = 16'h4353;
    tile_memory[ 61] = 16'hC7C7;
    tile_memory[ 62] = 16'h7FFF;
    tile_memory[ 63] = 16'h013D;
    tile_memory[ 64] = 16'h8585;
    tile_memory[ 65] = 16'h6724;
    tile_memory[ 66] = 16'hC3E3;
    tile_memory[ 67] = 16'hF7F1;
    tile_memory[ 68] = 16'hCFF7;
    tile_memory[ 69] = 16'h7FCF;
    tile_memory[ 70] = 16'hBE77;
    tile_memory[ 71] = 16'hE8AA;
    tile_memory[ 72] = 16'hF1D8;
    tile_memory[ 73] = 16'hFBFB;
    tile_memory[ 74] = 16'hB3FB;
    tile_memory[ 75] = 16'hF5B5;
    tile_memory[ 76] = 16'hEAE7;
    tile_memory[ 77] = 16'h2FAF;
    tile_memory[ 78] = 16'hA6A7;
    tile_memory[ 79] = 16'h7FBC;
    tile_memory[ 80] = 16'hDB7B;
    tile_memory[ 81] = 16'hC8DA;
    tile_memory[ 82] = 16'hF878;
    tile_memory[ 83] = 16'h8BF8;
    tile_memory[ 84] = 16'hFB3B;
    tile_memory[ 85] = 16'hF0F8;
    tile_memory[ 86] = 16'hDB9B;
    tile_memory[ 87] = 16'hF3DB;
    tile_memory[ 88] = 16'hEFFD;
    tile_memory[ 89] = 16'hF2FF;
    tile_memory[ 90] = 16'h4FB3;
    tile_memory[ 91] = 16'hDF5F;
    tile_memory[ 92] = 16'hC3D3;
    tile_memory[ 93] = 16'hC7C7;
    tile_memory[ 94] = 16'hFFFF;
    tile_memory[ 95] = 16'h01BD;
    tile_memory[ 96] = 16'h8787;
    tile_memory[ 97] = 16'h67A6;
    tile_memory[ 98] = 16'hC3E3;
    tile_memory[ 99] = 16'hF7F1;
    tile_memory[100] = 16'hEFF7;
    tile_memory[101] = 16'h7FEF;
    tile_memory[102] = 16'hBE77;
    tile_memory[103] = 16'hE9AA;
    tile_memory[104] = 16'hF9D9;
    tile_memory[105] = 16'hFBFB;
    tile_memory[106] = 16'hB3FB;
    tile_memory[107] = 16'hD5B5;
    tile_memory[108] = 16'hEAC7;
    tile_memory[109] = 16'hAFAF;
    tile_memory[110] = 16'hA6A7;
    tile_memory[111] = 16'h7FBC;
    tile_memory[112] = 16'hDF7F;
    tile_memory[113] = 16'hCCDA;
    tile_memory[114] = 16'hFC7C;
    tile_memory[115] = 16'h8BF8;
    tile_memory[116] = 16'hFB3B;
    tile_memory[117] = 16'hF2FA;
    tile_memory[118] = 16'hDB9B;
    tile_memory[119] = 16'hF3DB;
    tile_memory[120] = 16'hFFFD;
    tile_memory[121] = 16'hF6FF;
    tile_memory[122] = 16'h4FB7;
    tile_memory[123] = 16'hDF5F;
    tile_memory[124] = 16'hFBD3;
    tile_memory[125] = 16'hBFFF;
    tile_memory[126] = 16'h3FBF;
    tile_memory[127] = 16'h013D;
    tile_memory[128] = 16'h8787;
    tile_memory[129] = 16'h6766;
    tile_memory[130] = 16'hC3E3;
    tile_memory[131] = 16'hFDF9;
    tile_memory[132] = 16'hEDFD;
    tile_memory[133] = 16'h7FFF;
    tile_memory[134] = 16'h3E77;
    tile_memory[135] = 16'hE8AE;
    tile_memory[136] = 16'hF9D8;
    tile_memory[137] = 16'hFBFB;
    tile_memory[138] = 16'hB3FB;
    tile_memory[139] = 16'hF5B5;
    tile_memory[140] = 16'hEAE7;
    tile_memory[141] = 16'hAFAF;
    tile_memory[142] = 16'hA7A7;
    tile_memory[143] = 16'h7FBC;
    tile_memory[144] = 16'hDB7B;
    tile_memory[145] = 16'hDCDA;
    tile_memory[146] = 16'hFE7E;
    tile_memory[147] = 16'hCFFA;
    tile_memory[148] = 16'hFF3F;
    tile_memory[149] = 16'hF2FA;
    tile_memory[150] = 16'hDB9B;
    tile_memory[151] = 16'hF7DF;
    tile_memory[152] = 16'hEFFD;
    tile_memory[153] = 16'hF6FF;
    tile_memory[154] = 16'h4FF7;
    tile_memory[155] = 16'hDD5D;
    tile_memory[156] = 16'hFBDB;
    tile_memory[157] = 16'hB7FF;
    tile_memory[158] = 16'hBFBF;
    tile_memory[159] = 16'h01BD;
    tile_memory[160] = 16'hD797;
    tile_memory[161] = 16'h67E6;
    tile_memory[162] = 16'hC3E3;
    tile_memory[163] = 16'hFFF9;
    tile_memory[164] = 16'hEFFF;
    tile_memory[165] = 16'h7FFF;
    tile_memory[166] = 16'hBE77;
    tile_memory[167] = 16'hE9AA;
    tile_memory[168] = 16'hD9D9;
    tile_memory[169] = 16'hDBDB;
    tile_memory[170] = 16'hBBFB;
    tile_memory[171] = 16'hF5BD;
    tile_memory[172] = 16'hEEE7;
    tile_memory[173] = 16'hAFAF;
    tile_memory[174] = 16'hA7A7;
    tile_memory[175] = 16'h7FBC;
    tile_memory[176] = 16'hDF7B;
    tile_memory[177] = 16'hDDDF;
    tile_memory[178] = 16'hFF7F;
    tile_memory[179] = 16'h8FFB;
    tile_memory[180] = 16'hFF3F;
    tile_memory[181] = 16'hF2FE;
    tile_memory[182] = 16'hDB9B;
    tile_memory[183] = 16'hF7DF;
    tile_memory[184] = 16'hFFFD;
    tile_memory[185] = 16'hF6FF;
    tile_memory[186] = 16'hCFB7;
    tile_memory[187] = 16'hDFDF;
    tile_memory[188] = 16'hFBDB;
    tile_memory[189] = 16'hFFFF;
    tile_memory[190] = 16'hFFFF;
    tile_memory[191] = 16'h01FD;
    tile_memory[192] = 16'hC787;
    tile_memory[193] = 16'h67E6;
    tile_memory[194] = 16'hDBEB;
    tile_memory[195] = 16'hFDF9;
    tile_memory[196] = 16'hEDFD;
    tile_memory[197] = 16'h7FFF;
    tile_memory[198] = 16'h3E77;
    tile_memory[199] = 16'hEDAA;
    tile_memory[200] = 16'hFFDD;
    tile_memory[201] = 16'hFBFB;
    tile_memory[202] = 16'hBFFB;
    tile_memory[203] = 16'hF5BD;
    tile_memory[204] = 16'hEEE7;
    tile_memory[205] = 16'hAFAF;
    tile_memory[206] = 16'hA7A7;
    tile_memory[207] = 16'h7FBE;
    tile_memory[208] = 16'hDF7B;
    tile_memory[209] = 16'hDDDF;
    tile_memory[210] = 16'hFF7F;
    tile_memory[211] = 16'hCFFB;
    tile_memory[212] = 16'hFF3F;
    tile_memory[213] = 16'hF6FE;
    tile_memory[214] = 16'hDF9F;
    tile_memory[215] = 16'hF7DF;
    tile_memory[216] = 16'hEFFD;
    tile_memory[217] = 16'hF2FF;
    tile_memory[218] = 16'hDFB3;
    tile_memory[219] = 16'hDFDF;
    tile_memory[220] = 16'hFBDB;
    tile_memory[221] = 16'hFFFF;
    tile_memory[222] = 16'hFFFF;
    tile_memory[223] = 16'h01FF;
    tile_memory[224] = 16'h8787;
    tile_memory[225] = 16'h6FEF;
    tile_memory[226] = 16'hDBEB;
    tile_memory[227] = 16'hFFF9;
    tile_memory[228] = 16'hEFFF;
    tile_memory[229] = 16'h7FFF;
    tile_memory[230] = 16'hBE77;
    tile_memory[231] = 16'hEDAA;
    tile_memory[232] = 16'hFFDD;
    tile_memory[233] = 16'hFBFB;
    tile_memory[234] = 16'hBFFB;
    tile_memory[235] = 16'hF7BF;
    tile_memory[236] = 16'hEFFF;
    tile_memory[237] = 16'hAFAF;
    tile_memory[238] = 16'hB7B7;
    tile_memory[239] = 16'h7FBE;
    tile_memory[240] = 16'hFF7F;
    tile_memory[241] = 16'hCDDF;
    tile_memory[242] = 16'hFB7B;
    tile_memory[243] = 16'hCFFB;
    tile_memory[244] = 16'hFF3F;
    tile_memory[245] = 16'hF6FE;
    tile_memory[246] = 16'hDFBF;
    tile_memory[247] = 16'hF7DF;
    tile_memory[248] = 16'hFFFD;
    tile_memory[249] = 16'hF3FF;
    tile_memory[250] = 16'hCFF3;
    tile_memory[251] = 16'hDDDD;
    tile_memory[252] = 16'hFBDB;
    tile_memory[253] = 16'hFFFF;
    tile_memory[254] = 16'hFFFF;
    tile_memory[255] = 16'h01FF;
  end

endmodule
