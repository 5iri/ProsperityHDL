// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_1_enc_9_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h5AA0;
    tile_memory[  1] = 16'h69FE;
    tile_memory[  2] = 16'hDFFF;
    tile_memory[  3] = 16'hFF79;
    tile_memory[  4] = 16'h8FFF;
    tile_memory[  5] = 16'hFBB9;
    tile_memory[  6] = 16'hDAD9;
    tile_memory[  7] = 16'hFFB7;
    tile_memory[  8] = 16'hE971;
    tile_memory[  9] = 16'hFBF5;
    tile_memory[ 10] = 16'h48F7;
    tile_memory[ 11] = 16'hCFBB;
    tile_memory[ 12] = 16'h3FF7;
    tile_memory[ 13] = 16'hDF4C;
    tile_memory[ 14] = 16'h6FD3;
    tile_memory[ 15] = 16'hF6E0;
    tile_memory[ 16] = 16'hFF1A;
    tile_memory[ 17] = 16'h23B5;
    tile_memory[ 18] = 16'hF29E;
    tile_memory[ 19] = 16'hF6F3;
    tile_memory[ 20] = 16'h1EEB;
    tile_memory[ 21] = 16'hD7DE;
    tile_memory[ 22] = 16'h7F8E;
    tile_memory[ 23] = 16'hFE7D;
    tile_memory[ 24] = 16'hCF5D;
    tile_memory[ 25] = 16'hDFC2;
    tile_memory[ 26] = 16'h3D13;
    tile_memory[ 27] = 16'h0BFB;
    tile_memory[ 28] = 16'h7FFF;
    tile_memory[ 29] = 16'hB7AF;
    tile_memory[ 30] = 16'hBD5D;
    tile_memory[ 31] = 16'hE17F;
    tile_memory[ 32] = 16'h62FA;
    tile_memory[ 33] = 16'hDCF9;
    tile_memory[ 34] = 16'h8955;
    tile_memory[ 35] = 16'hDE2F;
    tile_memory[ 36] = 16'h73FA;
    tile_memory[ 37] = 16'hA7AC;
    tile_memory[ 38] = 16'h67E7;
    tile_memory[ 39] = 16'hE76D;
    tile_memory[ 40] = 16'hBFD3;
    tile_memory[ 41] = 16'hDAB9;
    tile_memory[ 42] = 16'hEB8B;
    tile_memory[ 43] = 16'hDD29;
    tile_memory[ 44] = 16'hFBF0;
    tile_memory[ 45] = 16'h979C;
    tile_memory[ 46] = 16'h7F77;
    tile_memory[ 47] = 16'hAEBF;
    tile_memory[ 48] = 16'h5AF4;
    tile_memory[ 49] = 16'hF7E6;
    tile_memory[ 50] = 16'hFD77;
    tile_memory[ 51] = 16'h7F5A;
    tile_memory[ 52] = 16'h976E;
    tile_memory[ 53] = 16'hFBF1;
    tile_memory[ 54] = 16'hDBCB;
    tile_memory[ 55] = 16'hFF8B;
    tile_memory[ 56] = 16'hC9CB;
    tile_memory[ 57] = 16'hE7E5;
    tile_memory[ 58] = 16'h2DD6;
    tile_memory[ 59] = 16'h671B;
    tile_memory[ 60] = 16'hAFBB;
    tile_memory[ 61] = 16'h97CC;
    tile_memory[ 62] = 16'hAC59;
    tile_memory[ 63] = 16'hE566;
    tile_memory[ 64] = 16'hE71C;
    tile_memory[ 65] = 16'h46D3;
    tile_memory[ 66] = 16'hF9DB;
    tile_memory[ 67] = 16'hD472;
    tile_memory[ 68] = 16'h2FEA;
    tile_memory[ 69] = 16'hDBDC;
    tile_memory[ 70] = 16'h7F8E;
    tile_memory[ 71] = 16'hD4F3;
    tile_memory[ 72] = 16'hDFAC;
    tile_memory[ 73] = 16'hD793;
    tile_memory[ 74] = 16'h7F12;
    tile_memory[ 75] = 16'h33FF;
    tile_memory[ 76] = 16'hFBEF;
    tile_memory[ 77] = 16'hA93B;
    tile_memory[ 78] = 16'hBF7F;
    tile_memory[ 79] = 16'hE8EF;
    tile_memory[ 80] = 16'h6FB2;
    tile_memory[ 81] = 16'hEFF8;
    tile_memory[ 82] = 16'hECD7;
    tile_memory[ 83] = 16'hCF15;
    tile_memory[ 84] = 16'h72F2;
    tile_memory[ 85] = 16'hF3B8;
    tile_memory[ 86] = 16'hADEF;
    tile_memory[ 87] = 16'hEF1D;
    tile_memory[ 88] = 16'hAFAF;
    tile_memory[ 89] = 16'h9BAB;
    tile_memory[ 90] = 16'hB38F;
    tile_memory[ 91] = 16'h7B3F;
    tile_memory[ 92] = 16'hDBB8;
    tile_memory[ 93] = 16'hEEBD;
    tile_memory[ 94] = 16'h7E3B;
    tile_memory[ 95] = 16'hEEBF;
    tile_memory[ 96] = 16'hFAC2;
    tile_memory[ 97] = 16'h5BFE;
    tile_memory[ 98] = 16'hDF1D;
    tile_memory[ 99] = 16'hFFFF;
    tile_memory[100] = 16'hBD6F;
    tile_memory[101] = 16'hFBB7;
    tile_memory[102] = 16'hFADB;
    tile_memory[103] = 16'hD74B;
    tile_memory[104] = 16'hEBF9;
    tile_memory[105] = 16'hF3AF;
    tile_memory[106] = 16'hF8F3;
    tile_memory[107] = 16'h8F3B;
    tile_memory[108] = 16'h7F3F;
    tile_memory[109] = 16'hA68E;
    tile_memory[110] = 16'hED15;
    tile_memory[111] = 16'hF6F9;
    tile_memory[112] = 16'h579D;
    tile_memory[113] = 16'h64F3;
    tile_memory[114] = 16'h3BFA;
    tile_memory[115] = 16'hF776;
    tile_memory[116] = 16'h0DFB;
    tile_memory[117] = 16'hC6FC;
    tile_memory[118] = 16'hFEBE;
    tile_memory[119] = 16'hF17E;
    tile_memory[120] = 16'hE776;
    tile_memory[121] = 16'hDFD7;
    tile_memory[122] = 16'hED10;
    tile_memory[123] = 16'h3AF1;
    tile_memory[124] = 16'hFBFD;
    tile_memory[125] = 16'hEBE7;
    tile_memory[126] = 16'hBFFD;
    tile_memory[127] = 16'hC77F;
    tile_memory[128] = 16'hFFDE;
    tile_memory[129] = 16'hFEF8;
    tile_memory[130] = 16'hBA4D;
    tile_memory[131] = 16'hFF74;
    tile_memory[132] = 16'h77F3;
    tile_memory[133] = 16'hABAE;
    tile_memory[134] = 16'hF5E7;
    tile_memory[135] = 16'hFFDE;
    tile_memory[136] = 16'hEFAD;
    tile_memory[137] = 16'hDCFB;
    tile_memory[138] = 16'h2FCA;
    tile_memory[139] = 16'hFB3F;
    tile_memory[140] = 16'hFBBF;
    tile_memory[141] = 16'hD6FF;
    tile_memory[142] = 16'h757C;
    tile_memory[143] = 16'hAFE7;
    tile_memory[144] = 16'h7FE0;
    tile_memory[145] = 16'hFD86;
    tile_memory[146] = 16'hDF3D;
    tile_memory[147] = 16'h7D5A;
    tile_memory[148] = 16'hFDE7;
    tile_memory[149] = 16'hFBE4;
    tile_memory[150] = 16'hDFFF;
    tile_memory[151] = 16'hE7D3;
    tile_memory[152] = 16'hFF28;
    tile_memory[153] = 16'hEA3F;
    tile_memory[154] = 16'hD9CE;
    tile_memory[155] = 16'h17BB;
    tile_memory[156] = 16'h3D75;
    tile_memory[157] = 16'hA44F;
    tile_memory[158] = 16'h4F79;
    tile_memory[159] = 16'hE3FB;
    tile_memory[160] = 16'h3DFD;
    tile_memory[161] = 16'h21F5;
    tile_memory[162] = 16'h319E;
    tile_memory[163] = 16'hDD7A;
    tile_memory[164] = 16'h6DEA;
    tile_memory[165] = 16'hF5FA;
    tile_memory[166] = 16'h7CED;
    tile_memory[167] = 16'hDBF5;
    tile_memory[168] = 16'hC7E4;
    tile_memory[169] = 16'h5EDA;
    tile_memory[170] = 16'h6F13;
    tile_memory[171] = 16'hA2EB;
    tile_memory[172] = 16'h7FFD;
    tile_memory[173] = 16'hB54B;
    tile_memory[174] = 16'hBD7F;
    tile_memory[175] = 16'hFB63;
    tile_memory[176] = 16'h56D7;
    tile_memory[177] = 16'hDEFA;
    tile_memory[178] = 16'hB37F;
    tile_memory[179] = 16'h7F66;
    tile_memory[180] = 16'hFB7A;
    tile_memory[181] = 16'hF7BA;
    tile_memory[182] = 16'hFD77;
    tile_memory[183] = 16'hDB4F;
    tile_memory[184] = 16'hFF55;
    tile_memory[185] = 16'h9EE9;
    tile_memory[186] = 16'hF38B;
    tile_memory[187] = 16'hDB69;
    tile_memory[188] = 16'hFFFD;
    tile_memory[189] = 16'h17DC;
    tile_memory[190] = 16'h3DD0;
    tile_memory[191] = 16'h6FAF;
    tile_memory[192] = 16'hFA8B;
    tile_memory[193] = 16'hC8DF;
    tile_memory[194] = 16'h8FDD;
    tile_memory[195] = 16'hDDF4;
    tile_memory[196] = 16'hFFEF;
    tile_memory[197] = 16'h7BFA;
    tile_memory[198] = 16'hFB5D;
    tile_memory[199] = 16'h478B;
    tile_memory[200] = 16'h5B3E;
    tile_memory[201] = 16'hF2ED;
    tile_memory[202] = 16'hA9DF;
    tile_memory[203] = 16'hAF1F;
    tile_memory[204] = 16'h357F;
    tile_memory[205] = 16'hD6BE;
    tile_memory[206] = 16'h1EB3;
    tile_memory[207] = 16'hE8E3;
    tile_memory[208] = 16'hEF5C;
    tile_memory[209] = 16'h2C99;
    tile_memory[210] = 16'hB3FB;
    tile_memory[211] = 16'hDBFB;
    tile_memory[212] = 16'hCFFE;
    tile_memory[213] = 16'hEBFC;
    tile_memory[214] = 16'h7FBC;
    tile_memory[215] = 16'hD9F3;
    tile_memory[216] = 16'hF77D;
    tile_memory[217] = 16'hF7A7;
    tile_memory[218] = 16'h79F1;
    tile_memory[219] = 16'hEBF9;
    tile_memory[220] = 16'h3B7D;
    tile_memory[221] = 16'hF953;
    tile_memory[222] = 16'hBD5D;
    tile_memory[223] = 16'hE4F7;
    tile_memory[224] = 16'h4EF2;
    tile_memory[225] = 16'hEFFF;
    tile_memory[226] = 16'h95EB;
    tile_memory[227] = 16'h2E6F;
    tile_memory[228] = 16'h7F77;
    tile_memory[229] = 16'hFBFB;
    tile_memory[230] = 16'hF5E5;
    tile_memory[231] = 16'hE75C;
    tile_memory[232] = 16'hEFF1;
    tile_memory[233] = 16'hB8BD;
    tile_memory[234] = 16'hE7EB;
    tile_memory[235] = 16'h57BF;
    tile_memory[236] = 16'hBEB8;
    tile_memory[237] = 16'h1EFC;
    tile_memory[238] = 16'h7DC1;
    tile_memory[239] = 16'hEE57;
    tile_memory[240] = 16'h5AC0;
    tile_memory[241] = 16'h41CE;
    tile_memory[242] = 16'hDF3D;
    tile_memory[243] = 16'hDF5E;
    tile_memory[244] = 16'hB566;
    tile_memory[245] = 16'h7BFB;
    tile_memory[246] = 16'hFACB;
    tile_memory[247] = 16'h4713;
    tile_memory[248] = 16'hE5A7;
    tile_memory[249] = 16'hFBA7;
    tile_memory[250] = 16'h28D5;
    tile_memory[251] = 16'h4F1B;
    tile_memory[252] = 16'h3DB7;
    tile_memory[253] = 16'hBC9D;
    tile_memory[254] = 16'hCC9D;
    tile_memory[255] = 16'hF761;
  end

endmodule
