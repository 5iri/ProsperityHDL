// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_1_enc_0_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h6100;
    tile_memory[  1] = 16'hAA00;
    tile_memory[  2] = 16'h0484;
    tile_memory[  3] = 16'h012D;
    tile_memory[  4] = 16'h41A9;
    tile_memory[  5] = 16'h0062;
    tile_memory[  6] = 16'h7130;
    tile_memory[  7] = 16'h4026;
    tile_memory[  8] = 16'h200B;
    tile_memory[  9] = 16'h0401;
    tile_memory[ 10] = 16'h4200;
    tile_memory[ 11] = 16'h3800;
    tile_memory[ 12] = 16'h3028;
    tile_memory[ 13] = 16'h404C;
    tile_memory[ 14] = 16'h0022;
    tile_memory[ 15] = 16'h1000;
    tile_memory[ 16] = 16'h1920;
    tile_memory[ 17] = 16'h3540;
    tile_memory[ 18] = 16'h1384;
    tile_memory[ 19] = 16'h8022;
    tile_memory[ 20] = 16'h84A4;
    tile_memory[ 21] = 16'h2002;
    tile_memory[ 22] = 16'h0020;
    tile_memory[ 23] = 16'h8421;
    tile_memory[ 24] = 16'h020D;
    tile_memory[ 25] = 16'h8880;
    tile_memory[ 26] = 16'h4100;
    tile_memory[ 27] = 16'h0A04;
    tile_memory[ 28] = 16'h6940;
    tile_memory[ 29] = 16'h4082;
    tile_memory[ 30] = 16'h2020;
    tile_memory[ 31] = 16'h0894;
    tile_memory[ 32] = 16'h2080;
    tile_memory[ 33] = 16'h20C8;
    tile_memory[ 34] = 16'h0140;
    tile_memory[ 35] = 16'h8944;
    tile_memory[ 36] = 16'h2004;
    tile_memory[ 37] = 16'h1440;
    tile_memory[ 38] = 16'h0369;
    tile_memory[ 39] = 16'h1140;
    tile_memory[ 40] = 16'h4440;
    tile_memory[ 41] = 16'h2208;
    tile_memory[ 42] = 16'hB351;
    tile_memory[ 43] = 16'h201E;
    tile_memory[ 44] = 16'h11C2;
    tile_memory[ 45] = 16'hA402;
    tile_memory[ 46] = 16'h7180;
    tile_memory[ 47] = 16'hC203;
    tile_memory[ 48] = 16'h8027;
    tile_memory[ 49] = 16'h0286;
    tile_memory[ 50] = 16'h1050;
    tile_memory[ 51] = 16'h1D40;
    tile_memory[ 52] = 16'h4045;
    tile_memory[ 53] = 16'h5030;
    tile_memory[ 54] = 16'h000A;
    tile_memory[ 55] = 16'h8090;
    tile_memory[ 56] = 16'h80A0;
    tile_memory[ 57] = 16'h0080;
    tile_memory[ 58] = 16'h001C;
    tile_memory[ 59] = 16'h1101;
    tile_memory[ 60] = 16'h0892;
    tile_memory[ 61] = 16'hE687;
    tile_memory[ 62] = 16'h0002;
    tile_memory[ 63] = 16'h208C;
    tile_memory[ 64] = 16'h0281;
    tile_memory[ 65] = 16'h2203;
    tile_memory[ 66] = 16'h8840;
    tile_memory[ 67] = 16'h01A0;
    tile_memory[ 68] = 16'h3246;
    tile_memory[ 69] = 16'h0840;
    tile_memory[ 70] = 16'hC800;
    tile_memory[ 71] = 16'h042A;
    tile_memory[ 72] = 16'h8200;
    tile_memory[ 73] = 16'h0042;
    tile_memory[ 74] = 16'h0090;
    tile_memory[ 75] = 16'h5540;
    tile_memory[ 76] = 16'h0201;
    tile_memory[ 77] = 16'h0A00;
    tile_memory[ 78] = 16'h0387;
    tile_memory[ 79] = 16'h3623;
    tile_memory[ 80] = 16'h8290;
    tile_memory[ 81] = 16'h0480;
    tile_memory[ 82] = 16'h4888;
    tile_memory[ 83] = 16'h8915;
    tile_memory[ 84] = 16'h0004;
    tile_memory[ 85] = 16'h0840;
    tile_memory[ 86] = 16'h21A0;
    tile_memory[ 87] = 16'h5412;
    tile_memory[ 88] = 16'h0804;
    tile_memory[ 89] = 16'h3003;
    tile_memory[ 90] = 16'h1028;
    tile_memory[ 91] = 16'hD01C;
    tile_memory[ 92] = 16'h2844;
    tile_memory[ 93] = 16'h8004;
    tile_memory[ 94] = 16'h2040;
    tile_memory[ 95] = 16'h0340;
    tile_memory[ 96] = 16'h05A0;
    tile_memory[ 97] = 16'h9050;
    tile_memory[ 98] = 16'h8863;
    tile_memory[ 99] = 16'h4C44;
    tile_memory[100] = 16'h5001;
    tile_memory[101] = 16'h4401;
    tile_memory[102] = 16'h3918;
    tile_memory[103] = 16'hC001;
    tile_memory[104] = 16'h0066;
    tile_memory[105] = 16'h2128;
    tile_memory[106] = 16'h0098;
    tile_memory[107] = 16'h7406;
    tile_memory[108] = 16'h0010;
    tile_memory[109] = 16'h0604;
    tile_memory[110] = 16'h2003;
    tile_memory[111] = 16'h0404;
    tile_memory[112] = 16'h0288;
    tile_memory[113] = 16'h0400;
    tile_memory[114] = 16'h1100;
    tile_memory[115] = 16'h00C8;
    tile_memory[116] = 16'h1642;
    tile_memory[117] = 16'h0444;
    tile_memory[118] = 16'h1000;
    tile_memory[119] = 16'h9900;
    tile_memory[120] = 16'h88A0;
    tile_memory[121] = 16'h1081;
    tile_memory[122] = 16'hF001;
    tile_memory[123] = 16'h0318;
    tile_memory[124] = 16'hA000;
    tile_memory[125] = 16'h0248;
    tile_memory[126] = 16'h1A06;
    tile_memory[127] = 16'h0240;
    tile_memory[128] = 16'h0014;
    tile_memory[129] = 16'hC4C0;
    tile_memory[130] = 16'h6AA4;
    tile_memory[131] = 16'h1404;
    tile_memory[132] = 16'h1844;
    tile_memory[133] = 16'h0040;
    tile_memory[134] = 16'h8020;
    tile_memory[135] = 16'h0011;
    tile_memory[136] = 16'h4034;
    tile_memory[137] = 16'h0C00;
    tile_memory[138] = 16'h0788;
    tile_memory[139] = 16'h1814;
    tile_memory[140] = 16'h1005;
    tile_memory[141] = 16'h8500;
    tile_memory[142] = 16'h0104;
    tile_memory[143] = 16'h0044;
    tile_memory[144] = 16'h3229;
    tile_memory[145] = 16'h0100;
    tile_memory[146] = 16'h1A62;
    tile_memory[147] = 16'h2C04;
    tile_memory[148] = 16'h58B0;
    tile_memory[149] = 16'hCC04;
    tile_memory[150] = 16'h1710;
    tile_memory[151] = 16'h1402;
    tile_memory[152] = 16'h09CE;
    tile_memory[153] = 16'h0200;
    tile_memory[154] = 16'h8008;
    tile_memory[155] = 16'h5292;
    tile_memory[156] = 16'h8500;
    tile_memory[157] = 16'h2300;
    tile_memory[158] = 16'h0008;
    tile_memory[159] = 16'h4500;
    tile_memory[160] = 16'h0200;
    tile_memory[161] = 16'h8061;
    tile_memory[162] = 16'h1204;
    tile_memory[163] = 16'h0302;
    tile_memory[164] = 16'h1150;
    tile_memory[165] = 16'h20C4;
    tile_memory[166] = 16'h08A0;
    tile_memory[167] = 16'h9000;
    tile_memory[168] = 16'h2102;
    tile_memory[169] = 16'h0122;
    tile_memory[170] = 16'h5000;
    tile_memory[171] = 16'h0104;
    tile_memory[172] = 16'hA881;
    tile_memory[173] = 16'hC058;
    tile_memory[174] = 16'h0288;
    tile_memory[175] = 16'h8052;
    tile_memory[176] = 16'h0010;
    tile_memory[177] = 16'h0001;
    tile_memory[178] = 16'h4081;
    tile_memory[179] = 16'h2000;
    tile_memory[180] = 16'h040C;
    tile_memory[181] = 16'h0102;
    tile_memory[182] = 16'h80A3;
    tile_memory[183] = 16'hD091;
    tile_memory[184] = 16'h0040;
    tile_memory[185] = 16'h0A40;
    tile_memory[186] = 16'h2004;
    tile_memory[187] = 16'h5074;
    tile_memory[188] = 16'h2000;
    tile_memory[189] = 16'h0011;
    tile_memory[190] = 16'h3010;
    tile_memory[191] = 16'h0100;
    tile_memory[192] = 16'h1008;
    tile_memory[193] = 16'h0014;
    tile_memory[194] = 16'h1002;
    tile_memory[195] = 16'h1800;
    tile_memory[196] = 16'h5020;
    tile_memory[197] = 16'hA000;
    tile_memory[198] = 16'h012A;
    tile_memory[199] = 16'h0400;
    tile_memory[200] = 16'h4064;
    tile_memory[201] = 16'h0084;
    tile_memory[202] = 16'h4040;
    tile_memory[203] = 16'h1A02;
    tile_memory[204] = 16'h1102;
    tile_memory[205] = 16'h0001;
    tile_memory[206] = 16'h2248;
    tile_memory[207] = 16'h3100;
    tile_memory[208] = 16'h8410;
    tile_memory[209] = 16'hC010;
    tile_memory[210] = 16'h1104;
    tile_memory[211] = 16'h0010;
    tile_memory[212] = 16'h1011;
    tile_memory[213] = 16'h2020;
    tile_memory[214] = 16'h0405;
    tile_memory[215] = 16'hC901;
    tile_memory[216] = 16'h1000;
    tile_memory[217] = 16'h0090;
    tile_memory[218] = 16'h8240;
    tile_memory[219] = 16'h0006;
    tile_memory[220] = 16'h90A0;
    tile_memory[221] = 16'h0040;
    tile_memory[222] = 16'h5A28;
    tile_memory[223] = 16'h4010;
    tile_memory[224] = 16'h0010;
    tile_memory[225] = 16'h0048;
    tile_memory[226] = 16'h684F;
    tile_memory[227] = 16'h0010;
    tile_memory[228] = 16'h0026;
    tile_memory[229] = 16'h0300;
    tile_memory[230] = 16'hA060;
    tile_memory[231] = 16'h8430;
    tile_memory[232] = 16'h4E04;
    tile_memory[233] = 16'h0224;
    tile_memory[234] = 16'h0011;
    tile_memory[235] = 16'h6094;
    tile_memory[236] = 16'h0040;
    tile_memory[237] = 16'h0110;
    tile_memory[238] = 16'h9010;
    tile_memory[239] = 16'h1120;
    tile_memory[240] = 16'h0528;
    tile_memory[241] = 16'h3004;
    tile_memory[242] = 16'h0202;
    tile_memory[243] = 16'h8408;
    tile_memory[244] = 16'h580C;
    tile_memory[245] = 16'h4908;
    tile_memory[246] = 16'h1010;
    tile_memory[247] = 16'h1204;
    tile_memory[248] = 16'h01C8;
    tile_memory[249] = 16'h5200;
    tile_memory[250] = 16'h0024;
    tile_memory[251] = 16'h1880;
    tile_memory[252] = 16'h2010;
    tile_memory[253] = 16'h0080;
    tile_memory[254] = 16'h0024;
    tile_memory[255] = 16'h7454;
  end

endmodule
