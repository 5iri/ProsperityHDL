// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_1_enc_2_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h1220;
    tile_memory[  1] = 16'h69FE;
    tile_memory[  2] = 16'h57FF;
    tile_memory[  3] = 16'hBB69;
    tile_memory[  4] = 16'h8F9F;
    tile_memory[  5] = 16'hBB39;
    tile_memory[  6] = 16'hD2D1;
    tile_memory[  7] = 16'hFDB4;
    tile_memory[  8] = 16'hA971;
    tile_memory[  9] = 16'hDBF5;
    tile_memory[ 10] = 16'h4077;
    tile_memory[ 11] = 16'hCFAB;
    tile_memory[ 12] = 16'h3BE7;
    tile_memory[ 13] = 16'hDB4C;
    tile_memory[ 14] = 16'h6FD3;
    tile_memory[ 15] = 16'hB6E0;
    tile_memory[ 16] = 16'hFF0A;
    tile_memory[ 17] = 16'h2335;
    tile_memory[ 18] = 16'hE294;
    tile_memory[ 19] = 16'hE6F1;
    tile_memory[ 20] = 16'h1EAB;
    tile_memory[ 21] = 16'hD7DE;
    tile_memory[ 22] = 16'h4F06;
    tile_memory[ 23] = 16'hBE3D;
    tile_memory[ 24] = 16'h4C5D;
    tile_memory[ 25] = 16'hCF42;
    tile_memory[ 26] = 16'h3C13;
    tile_memory[ 27] = 16'h09FB;
    tile_memory[ 28] = 16'h4DDB;
    tile_memory[ 29] = 16'h37AF;
    tile_memory[ 30] = 16'hB149;
    tile_memory[ 31] = 16'h213D;
    tile_memory[ 32] = 16'h60FA;
    tile_memory[ 33] = 16'hD459;
    tile_memory[ 34] = 16'h8954;
    tile_memory[ 35] = 16'hD20F;
    tile_memory[ 36] = 16'h41E8;
    tile_memory[ 37] = 16'hA7A4;
    tile_memory[ 38] = 16'h67C3;
    tile_memory[ 39] = 16'h6569;
    tile_memory[ 40] = 16'hB8D2;
    tile_memory[ 41] = 16'hCAB9;
    tile_memory[ 42] = 16'hCB83;
    tile_memory[ 43] = 16'hDC29;
    tile_memory[ 44] = 16'hF950;
    tile_memory[ 45] = 16'h939C;
    tile_memory[ 46] = 16'h5F77;
    tile_memory[ 47] = 16'h8EB9;
    tile_memory[ 48] = 16'h1874;
    tile_memory[ 49] = 16'hF7E6;
    tile_memory[ 50] = 16'h7567;
    tile_memory[ 51] = 16'h7B4A;
    tile_memory[ 52] = 16'h930E;
    tile_memory[ 53] = 16'hFBD1;
    tile_memory[ 54] = 16'hD1C3;
    tile_memory[ 55] = 16'hFD89;
    tile_memory[ 56] = 16'hC9CB;
    tile_memory[ 57] = 16'hC7E5;
    tile_memory[ 58] = 16'h2556;
    tile_memory[ 59] = 16'h6713;
    tile_memory[ 60] = 16'hAABB;
    tile_memory[ 61] = 16'h93CC;
    tile_memory[ 62] = 16'hA859;
    tile_memory[ 63] = 16'h2546;
    tile_memory[ 64] = 16'hE60C;
    tile_memory[ 65] = 16'h4653;
    tile_memory[ 66] = 16'hF9C3;
    tile_memory[ 67] = 16'hD420;
    tile_memory[ 68] = 16'h27A8;
    tile_memory[ 69] = 16'h5BDC;
    tile_memory[ 70] = 16'h6F0A;
    tile_memory[ 71] = 16'h84B3;
    tile_memory[ 72] = 16'hDEAC;
    tile_memory[ 73] = 16'hC713;
    tile_memory[ 74] = 16'h7E12;
    tile_memory[ 75] = 16'h317F;
    tile_memory[ 76] = 16'hD88B;
    tile_memory[ 77] = 16'h293B;
    tile_memory[ 78] = 16'h3B3A;
    tile_memory[ 79] = 16'hA8AD;
    tile_memory[ 80] = 16'h6D32;
    tile_memory[ 81] = 16'hEF58;
    tile_memory[ 82] = 16'hEC96;
    tile_memory[ 83] = 16'hC315;
    tile_memory[ 84] = 16'h40A0;
    tile_memory[ 85] = 16'hF3B0;
    tile_memory[ 86] = 16'hACCF;
    tile_memory[ 87] = 16'hEF19;
    tile_memory[ 88] = 16'h8AAE;
    tile_memory[ 89] = 16'h9B2B;
    tile_memory[ 90] = 16'h9385;
    tile_memory[ 91] = 16'h3A3F;
    tile_memory[ 92] = 16'hD998;
    tile_memory[ 93] = 16'hEEBD;
    tile_memory[ 94] = 16'h5E3B;
    tile_memory[ 95] = 16'hCABD;
    tile_memory[ 96] = 16'hB2C2;
    tile_memory[ 97] = 16'h5BFE;
    tile_memory[ 98] = 16'h4F09;
    tile_memory[ 99] = 16'hFFFF;
    tile_memory[100] = 16'hB96F;
    tile_memory[101] = 16'hBBB7;
    tile_memory[102] = 16'hF293;
    tile_memory[103] = 16'hD549;
    tile_memory[104] = 16'hEBF9;
    tile_memory[105] = 16'h93AF;
    tile_memory[106] = 16'hF873;
    tile_memory[107] = 16'h8F3B;
    tile_memory[108] = 16'h7B2F;
    tile_memory[109] = 16'hA28A;
    tile_memory[110] = 16'hED15;
    tile_memory[111] = 16'hB6D9;
    tile_memory[112] = 16'h578D;
    tile_memory[113] = 16'h64F3;
    tile_memory[114] = 16'h2BF0;
    tile_memory[115] = 16'hF736;
    tile_memory[116] = 16'h0DF9;
    tile_memory[117] = 16'h46FC;
    tile_memory[118] = 16'hEEB6;
    tile_memory[119] = 16'hB17E;
    tile_memory[120] = 16'hE676;
    tile_memory[121] = 16'hCF57;
    tile_memory[122] = 16'hE410;
    tile_memory[123] = 16'h3851;
    tile_memory[124] = 16'hDBED;
    tile_memory[125] = 16'hEBE7;
    tile_memory[126] = 16'h37E1;
    tile_memory[127] = 16'h877D;
    tile_memory[128] = 16'hFD5E;
    tile_memory[129] = 16'hFE78;
    tile_memory[130] = 16'hBA4D;
    tile_memory[131] = 16'hD374;
    tile_memory[132] = 16'h77B3;
    tile_memory[133] = 16'hA9A6;
    tile_memory[134] = 16'hF0E7;
    tile_memory[135] = 16'hFFDA;
    tile_memory[136] = 16'hCAAC;
    tile_memory[137] = 16'hDCFB;
    tile_memory[138] = 16'h2EC2;
    tile_memory[139] = 16'hF33F;
    tile_memory[140] = 16'hF99F;
    tile_memory[141] = 16'hD2FF;
    tile_memory[142] = 16'h717C;
    tile_memory[143] = 16'h8BE5;
    tile_memory[144] = 16'h35E0;
    tile_memory[145] = 16'hFD86;
    tile_memory[146] = 16'hDF39;
    tile_memory[147] = 16'h794A;
    tile_memory[148] = 16'hF8C5;
    tile_memory[149] = 16'hBBE4;
    tile_memory[150] = 16'hDDF7;
    tile_memory[151] = 16'hE7D2;
    tile_memory[152] = 16'hFF28;
    tile_memory[153] = 16'h8A1F;
    tile_memory[154] = 16'hD14E;
    tile_memory[155] = 16'h17A2;
    tile_memory[156] = 16'h3D75;
    tile_memory[157] = 16'hA04F;
    tile_memory[158] = 16'h4B79;
    tile_memory[159] = 16'h23DB;
    tile_memory[160] = 16'h3CFD;
    tile_memory[161] = 16'h21F5;
    tile_memory[162] = 16'h3194;
    tile_memory[163] = 16'h9D28;
    tile_memory[164] = 16'h6DEA;
    tile_memory[165] = 16'h757A;
    tile_memory[166] = 16'h7C69;
    tile_memory[167] = 16'hDBB5;
    tile_memory[168] = 16'h46E0;
    tile_memory[169] = 16'h5EDA;
    tile_memory[170] = 16'h6F13;
    tile_memory[171] = 16'hA26B;
    tile_memory[172] = 16'h6DAD;
    tile_memory[173] = 16'hB54B;
    tile_memory[174] = 16'h3C36;
    tile_memory[175] = 16'h3B61;
    tile_memory[176] = 16'h5657;
    tile_memory[177] = 16'h9ED2;
    tile_memory[178] = 16'hB33F;
    tile_memory[179] = 16'h5766;
    tile_memory[180] = 16'hC928;
    tile_memory[181] = 16'hF7B2;
    tile_memory[182] = 16'hFD53;
    tile_memory[183] = 16'hDB4F;
    tile_memory[184] = 16'hD854;
    tile_memory[185] = 16'h1EE9;
    tile_memory[186] = 16'hF301;
    tile_memory[187] = 16'h9B69;
    tile_memory[188] = 16'hFDFD;
    tile_memory[189] = 16'h13DC;
    tile_memory[190] = 16'h39D0;
    tile_memory[191] = 16'h6BAC;
    tile_memory[192] = 16'hF88B;
    tile_memory[193] = 16'hC8DB;
    tile_memory[194] = 16'h0FCD;
    tile_memory[195] = 16'h99E4;
    tile_memory[196] = 16'hFECF;
    tile_memory[197] = 16'h7B72;
    tile_memory[198] = 16'h795D;
    tile_memory[199] = 16'h478A;
    tile_memory[200] = 16'h1B3E;
    tile_memory[201] = 16'hF2ED;
    tile_memory[202] = 16'hA95F;
    tile_memory[203] = 16'hAE16;
    tile_memory[204] = 16'h356F;
    tile_memory[205] = 16'hD6BE;
    tile_memory[206] = 16'h1AB3;
    tile_memory[207] = 16'hE8E3;
    tile_memory[208] = 16'hEE5C;
    tile_memory[209] = 16'h2C99;
    tile_memory[210] = 16'hA3EB;
    tile_memory[211] = 16'h8BA9;
    tile_memory[212] = 16'hCFBC;
    tile_memory[213] = 16'h6BFC;
    tile_memory[214] = 16'h4F3C;
    tile_memory[215] = 16'h89B3;
    tile_memory[216] = 16'h7479;
    tile_memory[217] = 16'hA7A7;
    tile_memory[218] = 16'h78F1;
    tile_memory[219] = 16'hEB79;
    tile_memory[220] = 16'h083D;
    tile_memory[221] = 16'hF953;
    tile_memory[222] = 16'hBC18;
    tile_memory[223] = 16'h64B7;
    tile_memory[224] = 16'h4EF0;
    tile_memory[225] = 16'hEB5F;
    tile_memory[226] = 16'h95EA;
    tile_memory[227] = 16'h2E6F;
    tile_memory[228] = 16'h7D77;
    tile_memory[229] = 16'hFBF3;
    tile_memory[230] = 16'hF4C1;
    tile_memory[231] = 16'h6758;
    tile_memory[232] = 16'hECF0;
    tile_memory[233] = 16'h2835;
    tile_memory[234] = 16'hE7E1;
    tile_memory[235] = 16'h56BF;
    tile_memory[236] = 16'hB618;
    tile_memory[237] = 16'h1AEC;
    tile_memory[238] = 16'h5DC1;
    tile_memory[239] = 16'hCA53;
    tile_memory[240] = 16'h1240;
    tile_memory[241] = 16'h41CE;
    tile_memory[242] = 16'hDF3D;
    tile_memory[243] = 16'h9F5E;
    tile_memory[244] = 16'hB124;
    tile_memory[245] = 16'h7B7B;
    tile_memory[246] = 16'hF083;
    tile_memory[247] = 16'h4710;
    tile_memory[248] = 16'hE5A7;
    tile_memory[249] = 16'hBBA7;
    tile_memory[250] = 16'h2855;
    tile_memory[251] = 16'h4E1B;
    tile_memory[252] = 16'h39A7;
    tile_memory[253] = 16'hB89D;
    tile_memory[254] = 16'hCC9D;
    tile_memory[255] = 16'h3741;
  end

endmodule
