// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_v_enc_9_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h0004;
    tile_memory[  1] = 16'h6DEA;
    tile_memory[  2] = 16'h0270;
    tile_memory[  3] = 16'hEE78;
    tile_memory[  4] = 16'h8AF5;
    tile_memory[  5] = 16'h8202;
    tile_memory[  6] = 16'h2110;
    tile_memory[  7] = 16'h5CA2;
    tile_memory[  8] = 16'h2060;
    tile_memory[  9] = 16'h8931;
    tile_memory[ 10] = 16'h305E;
    tile_memory[ 11] = 16'h4802;
    tile_memory[ 12] = 16'h0F80;
    tile_memory[ 13] = 16'hCBA0;
    tile_memory[ 14] = 16'h2BD2;
    tile_memory[ 15] = 16'h5104;
    tile_memory[ 16] = 16'hED56;
    tile_memory[ 17] = 16'h280D;
    tile_memory[ 18] = 16'h6C8C;
    tile_memory[ 19] = 16'hD858;
    tile_memory[ 20] = 16'h98CB;
    tile_memory[ 21] = 16'h5190;
    tile_memory[ 22] = 16'h0002;
    tile_memory[ 23] = 16'h292A;
    tile_memory[ 24] = 16'h181F;
    tile_memory[ 25] = 16'hCC40;
    tile_memory[ 26] = 16'hF482;
    tile_memory[ 27] = 16'h4BEB;
    tile_memory[ 28] = 16'h4C26;
    tile_memory[ 29] = 16'h0723;
    tile_memory[ 30] = 16'h0C10;
    tile_memory[ 31] = 16'h8A0C;
    tile_memory[ 32] = 16'h02BE;
    tile_memory[ 33] = 16'h543B;
    tile_memory[ 34] = 16'h1124;
    tile_memory[ 35] = 16'h941C;
    tile_memory[ 36] = 16'h0880;
    tile_memory[ 37] = 16'h8C8C;
    tile_memory[ 38] = 16'hE267;
    tile_memory[ 39] = 16'h643D;
    tile_memory[ 40] = 16'h09F2;
    tile_memory[ 41] = 16'h4150;
    tile_memory[ 42] = 16'h8809;
    tile_memory[ 43] = 16'h0403;
    tile_memory[ 44] = 16'h0008;
    tile_memory[ 45] = 16'h73C4;
    tile_memory[ 46] = 16'h2339;
    tile_memory[ 47] = 16'h0948;
    tile_memory[ 48] = 16'h008D;
    tile_memory[ 49] = 16'h6DAA;
    tile_memory[ 50] = 16'h2222;
    tile_memory[ 51] = 16'hCA72;
    tile_memory[ 52] = 16'h87F0;
    tile_memory[ 53] = 16'hC882;
    tile_memory[ 54] = 16'hA140;
    tile_memory[ 55] = 16'h4CB1;
    tile_memory[ 56] = 16'h2600;
    tile_memory[ 57] = 16'h102D;
    tile_memory[ 58] = 16'hF444;
    tile_memory[ 59] = 16'h5020;
    tile_memory[ 60] = 16'h8D00;
    tile_memory[ 61] = 16'hC081;
    tile_memory[ 62] = 16'hA874;
    tile_memory[ 63] = 16'h4406;
    tile_memory[ 64] = 16'hE1D6;
    tile_memory[ 65] = 16'h6809;
    tile_memory[ 66] = 16'h7028;
    tile_memory[ 67] = 16'hB868;
    tile_memory[ 68] = 16'hA3DB;
    tile_memory[ 69] = 16'h4897;
    tile_memory[ 70] = 16'h8580;
    tile_memory[ 71] = 16'h1D02;
    tile_memory[ 72] = 16'hA80A;
    tile_memory[ 73] = 16'h0257;
    tile_memory[ 74] = 16'hE28A;
    tile_memory[ 75] = 16'h09A1;
    tile_memory[ 76] = 16'hCCAC;
    tile_memory[ 77] = 16'h118B;
    tile_memory[ 78] = 16'h6810;
    tile_memory[ 79] = 16'hAE00;
    tile_memory[ 80] = 16'h26BE;
    tile_memory[ 81] = 16'h857A;
    tile_memory[ 82] = 16'h1110;
    tile_memory[ 83] = 16'h8015;
    tile_memory[ 84] = 16'h24B0;
    tile_memory[ 85] = 16'h848D;
    tile_memory[ 86] = 16'h912F;
    tile_memory[ 87] = 16'hA43D;
    tile_memory[ 88] = 16'h3280;
    tile_memory[ 89] = 16'h2150;
    tile_memory[ 90] = 16'hC88A;
    tile_memory[ 91] = 16'h1803;
    tile_memory[ 92] = 16'h0208;
    tile_memory[ 93] = 16'h512C;
    tile_memory[ 94] = 16'h317C;
    tile_memory[ 95] = 16'h0C40;
    tile_memory[ 96] = 16'h0084;
    tile_memory[ 97] = 16'h6422;
    tile_memory[ 98] = 16'h0265;
    tile_memory[ 99] = 16'hCC58;
    tile_memory[100] = 16'h8EE0;
    tile_memory[101] = 16'h0802;
    tile_memory[102] = 16'h3340;
    tile_memory[103] = 16'h4AA2;
    tile_memory[104] = 16'h0EE8;
    tile_memory[105] = 16'h00BB;
    tile_memory[106] = 16'h324C;
    tile_memory[107] = 16'h4102;
    tile_memory[108] = 16'h0C01;
    tile_memory[109] = 16'h4081;
    tile_memory[110] = 16'hA890;
    tile_memory[111] = 16'h4000;
    tile_memory[112] = 16'hF1D4;
    tile_memory[113] = 16'h2489;
    tile_memory[114] = 16'h609C;
    tile_memory[115] = 16'h9808;
    tile_memory[116] = 16'hC0CB;
    tile_memory[117] = 16'h0893;
    tile_memory[118] = 16'h0400;
    tile_memory[119] = 16'h291B;
    tile_memory[120] = 16'h080E;
    tile_memory[121] = 16'h0040;
    tile_memory[122] = 16'hE022;
    tile_memory[123] = 16'hA92B;
    tile_memory[124] = 16'hC424;
    tile_memory[125] = 16'h2123;
    tile_memory[126] = 16'h0813;
    tile_memory[127] = 16'h2214;
    tile_memory[128] = 16'h46B8;
    tile_memory[129] = 16'hB431;
    tile_memory[130] = 16'h1580;
    tile_memory[131] = 16'h0152;
    tile_memory[132] = 16'h1C92;
    tile_memory[133] = 16'h0A68;
    tile_memory[134] = 16'h04AD;
    tile_memory[135] = 16'hA45F;
    tile_memory[136] = 16'h305C;
    tile_memory[137] = 16'h0951;
    tile_memory[138] = 16'h0888;
    tile_memory[139] = 16'h2493;
    tile_memory[140] = 16'h420B;
    tile_memory[141] = 16'h7702;
    tile_memory[142] = 16'h2138;
    tile_memory[143] = 16'hAC08;
    tile_memory[144] = 16'h0084;
    tile_memory[145] = 16'h7D2A;
    tile_memory[146] = 16'h002A;
    tile_memory[147] = 16'h4C50;
    tile_memory[148] = 16'h82E0;
    tile_memory[149] = 16'h6302;
    tile_memory[150] = 16'h2100;
    tile_memory[151] = 16'h4CA2;
    tile_memory[152] = 16'hC0C0;
    tile_memory[153] = 16'h0139;
    tile_memory[154] = 16'h704F;
    tile_memory[155] = 16'h0023;
    tile_memory[156] = 16'h0408;
    tile_memory[157] = 16'h4080;
    tile_memory[158] = 16'h0910;
    tile_memory[159] = 16'h4000;
    tile_memory[160] = 16'hF5D4;
    tile_memory[161] = 16'h6809;
    tile_memory[162] = 16'h408C;
    tile_memory[163] = 16'h9900;
    tile_memory[164] = 16'hA0CA;
    tile_memory[165] = 16'h0297;
    tile_memory[166] = 16'h2000;
    tile_memory[167] = 16'h290B;
    tile_memory[168] = 16'h080E;
    tile_memory[169] = 16'h0200;
    tile_memory[170] = 16'hE088;
    tile_memory[171] = 16'h4863;
    tile_memory[172] = 16'h5824;
    tile_memory[173] = 16'h0302;
    tile_memory[174] = 16'h0814;
    tile_memory[175] = 16'h2204;
    tile_memory[176] = 16'h46B4;
    tile_memory[177] = 16'h04E0;
    tile_memory[178] = 16'h1000;
    tile_memory[179] = 16'hC414;
    tile_memory[180] = 16'h1C80;
    tile_memory[181] = 16'h0DC8;
    tile_memory[182] = 16'h8067;
    tile_memory[183] = 16'h8E5D;
    tile_memory[184] = 16'h0290;
    tile_memory[185] = 16'h414A;
    tile_memory[186] = 16'h4CC8;
    tile_memory[187] = 16'h0453;
    tile_memory[188] = 16'h400B;
    tile_memory[189] = 16'h6820;
    tile_memory[190] = 16'h2128;
    tile_memory[191] = 16'h0948;
    tile_memory[192] = 16'h0084;
    tile_memory[193] = 16'h660A;
    tile_memory[194] = 16'h002A;
    tile_memory[195] = 16'h4C50;
    tile_memory[196] = 16'h8EE2;
    tile_memory[197] = 16'h8002;
    tile_memory[198] = 16'h3100;
    tile_memory[199] = 16'h40A2;
    tile_memory[200] = 16'h4000;
    tile_memory[201] = 16'h042D;
    tile_memory[202] = 16'hB24F;
    tile_memory[203] = 16'h1100;
    tile_memory[204] = 16'h0C08;
    tile_memory[205] = 16'hC080;
    tile_memory[206] = 16'h0812;
    tile_memory[207] = 16'h4001;
    tile_memory[208] = 16'hD154;
    tile_memory[209] = 16'h2089;
    tile_memory[210] = 16'h488C;
    tile_memory[211] = 16'h9888;
    tile_memory[212] = 16'hA0CE;
    tile_memory[213] = 16'h023A;
    tile_memory[214] = 16'h8000;
    tile_memory[215] = 16'h0902;
    tile_memory[216] = 16'h800E;
    tile_memory[217] = 16'h0200;
    tile_memory[218] = 16'hE08A;
    tile_memory[219] = 16'h6B61;
    tile_memory[220] = 16'h44A4;
    tile_memory[221] = 16'h2183;
    tile_memory[222] = 16'h0815;
    tile_memory[223] = 16'h0A10;
    tile_memory[224] = 16'h22A4;
    tile_memory[225] = 16'h4078;
    tile_memory[226] = 16'h1180;
    tile_memory[227] = 16'h8010;
    tile_memory[228] = 16'h0C00;
    tile_memory[229] = 16'h0E8A;
    tile_memory[230] = 16'h8047;
    tile_memory[231] = 16'h285D;
    tile_memory[232] = 16'h0210;
    tile_memory[233] = 16'h1150;
    tile_memory[234] = 16'hE888;
    tile_memory[235] = 16'h00D3;
    tile_memory[236] = 16'h0108;
    tile_memory[237] = 16'h6100;
    tile_memory[238] = 16'h6128;
    tile_memory[239] = 16'h8940;
    tile_memory[240] = 16'h0084;
    tile_memory[241] = 16'hE446;
    tile_memory[242] = 16'h00A2;
    tile_memory[243] = 16'h4D50;
    tile_memory[244] = 16'h8260;
    tile_memory[245] = 16'h2002;
    tile_memory[246] = 16'h2900;
    tile_memory[247] = 16'h3AA6;
    tile_memory[248] = 16'hC401;
    tile_memory[249] = 16'h00A5;
    tile_memory[250] = 16'h514F;
    tile_memory[251] = 16'h0202;
    tile_memory[252] = 16'h0418;
    tile_memory[253] = 16'h7080;
    tile_memory[254] = 16'h0850;
    tile_memory[255] = 16'h4206;
  end

endmodule
