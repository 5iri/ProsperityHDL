// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module attention_enc_1_q_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h4B30;
    tile_memory[  1] = 16'h672D;
    tile_memory[  2] = 16'h0340;
    tile_memory[  3] = 16'hBB20;
    tile_memory[  4] = 16'h100A;
    tile_memory[  5] = 16'h0014;
    tile_memory[  6] = 16'h0645;
    tile_memory[  7] = 16'h0200;
    tile_memory[  8] = 16'h0E01;
    tile_memory[  9] = 16'hE91C;
    tile_memory[ 10] = 16'h3C20;
    tile_memory[ 11] = 16'h0F40;
    tile_memory[ 12] = 16'hA780;
    tile_memory[ 13] = 16'hE023;
    tile_memory[ 14] = 16'h302E;
    tile_memory[ 15] = 16'h0080;
    tile_memory[ 16] = 16'h8800;
    tile_memory[ 17] = 16'hA400;
    tile_memory[ 18] = 16'h2812;
    tile_memory[ 19] = 16'h8852;
    tile_memory[ 20] = 16'h0018;
    tile_memory[ 21] = 16'h420A;
    tile_memory[ 22] = 16'h0516;
    tile_memory[ 23] = 16'h8355;
    tile_memory[ 24] = 16'h4330;
    tile_memory[ 25] = 16'h45A1;
    tile_memory[ 26] = 16'h0340;
    tile_memory[ 27] = 16'h936A;
    tile_memory[ 28] = 16'h1522;
    tile_memory[ 29] = 16'h8014;
    tile_memory[ 30] = 16'h0041;
    tile_memory[ 31] = 16'h2200;
    tile_memory[ 32] = 16'h4E01;
    tile_memory[ 33] = 16'hB108;
    tile_memory[ 34] = 16'h3828;
    tile_memory[ 35] = 16'h0E40;
    tile_memory[ 36] = 16'h0300;
    tile_memory[ 37] = 16'h0812;
    tile_memory[ 38] = 16'h22AC;
    tile_memory[ 39] = 16'h41A0;
    tile_memory[ 40] = 16'h0822;
    tile_memory[ 41] = 16'hA000;
    tile_memory[ 42] = 16'h2822;
    tile_memory[ 43] = 16'h8853;
    tile_memory[ 44] = 16'h4018;
    tile_memory[ 45] = 16'h9712;
    tile_memory[ 46] = 16'h0150;
    tile_memory[ 47] = 16'h4250;
    tile_memory[ 48] = 16'h4130;
    tile_memory[ 49] = 16'h4721;
    tile_memory[ 50] = 16'h0242;
    tile_memory[ 51] = 16'h5308;
    tile_memory[ 52] = 16'h1502;
    tile_memory[ 53] = 16'h8014;
    tile_memory[ 54] = 16'h88C0;
    tile_memory[ 55] = 16'h2240;
    tile_memory[ 56] = 16'h2A01;
    tile_memory[ 57] = 16'hA00A;
    tile_memory[ 58] = 16'hB828;
    tile_memory[ 59] = 16'h0628;
    tile_memory[ 60] = 16'h7B32;
    tile_memory[ 61] = 16'h6A32;
    tile_memory[ 62] = 16'h02AC;
    tile_memory[ 63] = 16'h0288;
    tile_memory[ 64] = 16'h0C60;
    tile_memory[ 65] = 16'hA048;
    tile_memory[ 66] = 16'h2832;
    tile_memory[ 67] = 16'h8853;
    tile_memory[ 68] = 16'h8418;
    tile_memory[ 69] = 16'h9230;
    tile_memory[ 70] = 16'h2140;
    tile_memory[ 71] = 16'h4211;
    tile_memory[ 72] = 16'h4230;
    tile_memory[ 73] = 16'hA500;
    tile_memory[ 74] = 16'h19E8;
    tile_memory[ 75] = 16'hF78A;
    tile_memory[ 76] = 16'h162A;
    tile_memory[ 77] = 16'h8010;
    tile_memory[ 78] = 16'h4460;
    tile_memory[ 79] = 16'h325C;
    tile_memory[ 80] = 16'h5242;
    tile_memory[ 81] = 16'h500C;
    tile_memory[ 82] = 16'hBC28;
    tile_memory[ 83] = 16'h0E60;
    tile_memory[ 84] = 16'hFF20;
    tile_memory[ 85] = 16'hF837;
    tile_memory[ 86] = 16'h362C;
    tile_memory[ 87] = 16'h26AA;
    tile_memory[ 88] = 16'h8C70;
    tile_memory[ 89] = 16'hA018;
    tile_memory[ 90] = 16'h3876;
    tile_memory[ 91] = 16'h0052;
    tile_memory[ 92] = 16'h8013;
    tile_memory[ 93] = 16'h8221;
    tile_memory[ 94] = 16'h6010;
    tile_memory[ 95] = 16'h4251;
    tile_memory[ 96] = 16'h0200;
    tile_memory[ 97] = 16'h6500;
    tile_memory[ 98] = 16'h0A62;
    tile_memory[ 99] = 16'hDBCA;
    tile_memory[100] = 16'h170A;
    tile_memory[101] = 16'h8010;
    tile_memory[102] = 16'h4860;
    tile_memory[103] = 16'h30B4;
    tile_memory[104] = 16'h4A40;
    tile_memory[105] = 16'h591C;
    tile_memory[106] = 16'hBC28;
    tile_memory[107] = 16'h0F48;
    tile_memory[108] = 16'hE624;
    tile_memory[109] = 16'h66B3;
    tile_memory[110] = 16'h242C;
    tile_memory[111] = 16'h0208;
    tile_memory[112] = 16'h0C30;
    tile_memory[113] = 16'hB000;
    tile_memory[114] = 16'h2022;
    tile_memory[115] = 16'hA252;
    tile_memory[116] = 16'h9421;
    tile_memory[117] = 16'h8210;
    tile_memory[118] = 16'h2418;
    tile_memory[119] = 16'h1115;
    tile_memory[120] = 16'h0101;
    tile_memory[121] = 16'h4500;
    tile_memory[122] = 16'h21C0;
    tile_memory[123] = 16'h3B28;
    tile_memory[124] = 16'h930A;
    tile_memory[125] = 16'h0010;
    tile_memory[126] = 16'h0861;
    tile_memory[127] = 16'h3060;
    tile_memory[128] = 16'h4A00;
    tile_memory[129] = 16'hC008;
    tile_memory[130] = 16'h35A8;
    tile_memory[131] = 16'h0B40;
    tile_memory[132] = 16'hE300;
    tile_memory[133] = 16'h2003;
    tile_memory[134] = 16'h3020;
    tile_memory[135] = 16'h6681;
    tile_memory[136] = 16'h8C40;
    tile_memory[137] = 16'h8000;
    tile_memory[138] = 16'hA000;
    tile_memory[139] = 16'h8858;
    tile_memory[140] = 16'h9419;
    tile_memory[141] = 16'h9512;
    tile_memory[142] = 16'h0108;
    tile_memory[143] = 16'h5101;
    tile_memory[144] = 16'h0201;
    tile_memory[145] = 16'h6580;
    tile_memory[146] = 16'h0240;
    tile_memory[147] = 16'hCD00;
    tile_memory[148] = 16'h1002;
    tile_memory[149] = 16'h0010;
    tile_memory[150] = 16'h0040;
    tile_memory[151] = 16'h0023;
    tile_memory[152] = 16'h42C2;
    tile_memory[153] = 16'h5988;
    tile_memory[154] = 16'h3828;
    tile_memory[155] = 16'h0A40;
    tile_memory[156] = 16'hA214;
    tile_memory[157] = 16'h2233;
    tile_memory[158] = 16'hA02C;
    tile_memory[159] = 16'h0201;
    tile_memory[160] = 16'h0C28;
    tile_memory[161] = 16'h9000;
    tile_memory[162] = 16'hA812;
    tile_memory[163] = 16'h8052;
    tile_memory[164] = 16'h9018;
    tile_memory[165] = 16'h0202;
    tile_memory[166] = 16'h2400;
    tile_memory[167] = 16'h4201;
    tile_memory[168] = 16'h0001;
    tile_memory[169] = 16'h6D84;
    tile_memory[170] = 16'h0A40;
    tile_memory[171] = 16'h8730;
    tile_memory[172] = 16'h1422;
    tile_memory[173] = 16'h8010;
    tile_memory[174] = 16'h0255;
    tile_memory[175] = 16'h3180;
    tile_memory[176] = 16'h4E80;
    tile_memory[177] = 16'h711D;
    tile_memory[178] = 16'h2C29;
    tile_memory[179] = 16'h8D41;
    tile_memory[180] = 16'h8310;
    tile_memory[181] = 16'h6433;
    tile_memory[182] = 16'hA028;
    tile_memory[183] = 16'h0F05;
    tile_memory[184] = 16'h0020;
    tile_memory[185] = 16'h8000;
    tile_memory[186] = 16'hAC02;
    tile_memory[187] = 16'h8092;
    tile_memory[188] = 16'h9412;
    tile_memory[189] = 16'hAA22;
    tile_memory[190] = 16'h0648;
    tile_memory[191] = 16'h4B57;
    tile_memory[192] = 16'h4203;
    tile_memory[193] = 16'h4500;
    tile_memory[194] = 16'h0B60;
    tile_memory[195] = 16'h9BB8;
    tile_memory[196] = 16'h970A;
    tile_memory[197] = 16'h9014;
    tile_memory[198] = 16'h0645;
    tile_memory[199] = 16'h118C;
    tile_memory[200] = 16'h5E11;
    tile_memory[201] = 16'hF91F;
    tile_memory[202] = 16'hBC29;
    tile_memory[203] = 16'h0B41;
    tile_memory[204] = 16'hA294;
    tile_memory[205] = 16'h7037;
    tile_memory[206] = 16'hE028;
    tile_memory[207] = 16'h6320;
    tile_memory[208] = 16'h2C30;
    tile_memory[209] = 16'h8000;
    tile_memory[210] = 16'hACB2;
    tile_memory[211] = 16'h8052;
    tile_memory[212] = 16'h9031;
    tile_memory[213] = 16'h8602;
    tile_memory[214] = 16'h4450;
    tile_memory[215] = 16'hCB51;
    tile_memory[216] = 16'h0121;
    tile_memory[217] = 16'h4500;
    tile_memory[218] = 16'h0940;
    tile_memory[219] = 16'h93C8;
    tile_memory[220] = 16'h8212;
    tile_memory[221] = 16'h9034;
    tile_memory[222] = 16'h0044;
    tile_memory[223] = 16'h30CC;
    tile_memory[224] = 16'h4620;
    tile_memory[225] = 16'hF11D;
    tile_memory[226] = 16'hBC01;
    tile_memory[227] = 16'h0B40;
    tile_memory[228] = 16'hA284;
    tile_memory[229] = 16'h7211;
    tile_memory[230] = 16'h0008;
    tile_memory[231] = 16'h2228;
    tile_memory[232] = 16'h0020;
    tile_memory[233] = 16'h2000;
    tile_memory[234] = 16'hB432;
    tile_memory[235] = 16'h80D0;
    tile_memory[236] = 16'h9014;
    tile_memory[237] = 16'h8622;
    tile_memory[238] = 16'h4408;
    tile_memory[239] = 16'hCB53;
    tile_memory[240] = 16'h0B21;
    tile_memory[241] = 16'h4504;
    tile_memory[242] = 16'h8140;
    tile_memory[243] = 16'h93C8;
    tile_memory[244] = 16'h924A;
    tile_memory[245] = 16'h0004;
    tile_memory[246] = 16'h0040;
    tile_memory[247] = 16'h3084;
    tile_memory[248] = 16'h4A00;
    tile_memory[249] = 16'h7008;
    tile_memory[250] = 16'hBCA8;
    tile_memory[251] = 16'h0B60;
    tile_memory[252] = 16'hE300;
    tile_memory[253] = 16'h6233;
    tile_memory[254] = 16'h0004;
    tile_memory[255] = 16'h2200;
  end

endmodule
