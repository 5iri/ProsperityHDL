// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module attention_enc_1_q_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h4B30;  // Neuron 0
    neuron_patterns[  1] = 16'h672D;  // Neuron 1
    neuron_patterns[  2] = 16'h0340;  // Neuron 2
    neuron_patterns[  3] = 16'hBB20;  // Neuron 3
    neuron_patterns[  4] = 16'h100A;  // Neuron 4
    neuron_patterns[  5] = 16'h0014;  // Neuron 5
    neuron_patterns[  6] = 16'h0645;  // Neuron 6
    neuron_patterns[  7] = 16'h0200;  // Neuron 7
    neuron_patterns[  8] = 16'h0E01;  // Neuron 8
    neuron_patterns[  9] = 16'hE91C;  // Neuron 9
    neuron_patterns[ 10] = 16'h3C20;  // Neuron 10
    neuron_patterns[ 11] = 16'h0F40;  // Neuron 11
    neuron_patterns[ 12] = 16'hA780;  // Neuron 12
    neuron_patterns[ 13] = 16'hE023;  // Neuron 13
    neuron_patterns[ 14] = 16'h302E;  // Neuron 14
    neuron_patterns[ 15] = 16'h0080;  // Neuron 15
    neuron_patterns[ 16] = 16'h8800;  // Neuron 16
    neuron_patterns[ 17] = 16'hA400;  // Neuron 17
    neuron_patterns[ 18] = 16'h2812;  // Neuron 18
    neuron_patterns[ 19] = 16'h8852;  // Neuron 19
    neuron_patterns[ 20] = 16'h0018;  // Neuron 20
    neuron_patterns[ 21] = 16'h420A;  // Neuron 21
    neuron_patterns[ 22] = 16'h0516;  // Neuron 22
    neuron_patterns[ 23] = 16'h8355;  // Neuron 23
    neuron_patterns[ 24] = 16'h4330;  // Neuron 24
    neuron_patterns[ 25] = 16'h45A1;  // Neuron 25
    neuron_patterns[ 26] = 16'h0340;  // Neuron 26
    neuron_patterns[ 27] = 16'h936A;  // Neuron 27
    neuron_patterns[ 28] = 16'h1522;  // Neuron 28
    neuron_patterns[ 29] = 16'h8014;  // Neuron 29
    neuron_patterns[ 30] = 16'h0041;  // Neuron 30
    neuron_patterns[ 31] = 16'h2200;  // Neuron 31
    neuron_patterns[ 32] = 16'h4E01;  // Neuron 32
    neuron_patterns[ 33] = 16'hB108;  // Neuron 33
    neuron_patterns[ 34] = 16'h3828;  // Neuron 34
    neuron_patterns[ 35] = 16'h0E40;  // Neuron 35
    neuron_patterns[ 36] = 16'h0300;  // Neuron 36
    neuron_patterns[ 37] = 16'h0812;  // Neuron 37
    neuron_patterns[ 38] = 16'h22AC;  // Neuron 38
    neuron_patterns[ 39] = 16'h41A0;  // Neuron 39
    neuron_patterns[ 40] = 16'h0822;  // Neuron 40
    neuron_patterns[ 41] = 16'hA000;  // Neuron 41
    neuron_patterns[ 42] = 16'h2822;  // Neuron 42
    neuron_patterns[ 43] = 16'h8853;  // Neuron 43
    neuron_patterns[ 44] = 16'h4018;  // Neuron 44
    neuron_patterns[ 45] = 16'h9712;  // Neuron 45
    neuron_patterns[ 46] = 16'h0150;  // Neuron 46
    neuron_patterns[ 47] = 16'h4250;  // Neuron 47
    neuron_patterns[ 48] = 16'h4130;  // Neuron 48
    neuron_patterns[ 49] = 16'h4721;  // Neuron 49
    neuron_patterns[ 50] = 16'h0242;  // Neuron 50
    neuron_patterns[ 51] = 16'h5308;  // Neuron 51
    neuron_patterns[ 52] = 16'h1502;  // Neuron 52
    neuron_patterns[ 53] = 16'h8014;  // Neuron 53
    neuron_patterns[ 54] = 16'h88C0;  // Neuron 54
    neuron_patterns[ 55] = 16'h2240;  // Neuron 55
    neuron_patterns[ 56] = 16'h2A01;  // Neuron 56
    neuron_patterns[ 57] = 16'hA00A;  // Neuron 57
    neuron_patterns[ 58] = 16'hB828;  // Neuron 58
    neuron_patterns[ 59] = 16'h0628;  // Neuron 59
    neuron_patterns[ 60] = 16'h7B32;  // Neuron 60
    neuron_patterns[ 61] = 16'h6A32;  // Neuron 61
    neuron_patterns[ 62] = 16'h02AC;  // Neuron 62
    neuron_patterns[ 63] = 16'h0288;  // Neuron 63
    neuron_patterns[ 64] = 16'h0C60;  // Neuron 64
    neuron_patterns[ 65] = 16'hA048;  // Neuron 65
    neuron_patterns[ 66] = 16'h2832;  // Neuron 66
    neuron_patterns[ 67] = 16'h8853;  // Neuron 67
    neuron_patterns[ 68] = 16'h8418;  // Neuron 68
    neuron_patterns[ 69] = 16'h9230;  // Neuron 69
    neuron_patterns[ 70] = 16'h2140;  // Neuron 70
    neuron_patterns[ 71] = 16'h4211;  // Neuron 71
    neuron_patterns[ 72] = 16'h4230;  // Neuron 72
    neuron_patterns[ 73] = 16'hA500;  // Neuron 73
    neuron_patterns[ 74] = 16'h19E8;  // Neuron 74
    neuron_patterns[ 75] = 16'hF78A;  // Neuron 75
    neuron_patterns[ 76] = 16'h162A;  // Neuron 76
    neuron_patterns[ 77] = 16'h8010;  // Neuron 77
    neuron_patterns[ 78] = 16'h4460;  // Neuron 78
    neuron_patterns[ 79] = 16'h325C;  // Neuron 79
    neuron_patterns[ 80] = 16'h5242;  // Neuron 80
    neuron_patterns[ 81] = 16'h500C;  // Neuron 81
    neuron_patterns[ 82] = 16'hBC28;  // Neuron 82
    neuron_patterns[ 83] = 16'h0E60;  // Neuron 83
    neuron_patterns[ 84] = 16'hFF20;  // Neuron 84
    neuron_patterns[ 85] = 16'hF837;  // Neuron 85
    neuron_patterns[ 86] = 16'h362C;  // Neuron 86
    neuron_patterns[ 87] = 16'h26AA;  // Neuron 87
    neuron_patterns[ 88] = 16'h8C70;  // Neuron 88
    neuron_patterns[ 89] = 16'hA018;  // Neuron 89
    neuron_patterns[ 90] = 16'h3876;  // Neuron 90
    neuron_patterns[ 91] = 16'h0052;  // Neuron 91
    neuron_patterns[ 92] = 16'h8013;  // Neuron 92
    neuron_patterns[ 93] = 16'h8221;  // Neuron 93
    neuron_patterns[ 94] = 16'h6010;  // Neuron 94
    neuron_patterns[ 95] = 16'h4251;  // Neuron 95
    neuron_patterns[ 96] = 16'h0200;  // Neuron 96
    neuron_patterns[ 97] = 16'h6500;  // Neuron 97
    neuron_patterns[ 98] = 16'h0A62;  // Neuron 98
    neuron_patterns[ 99] = 16'hDBCA;  // Neuron 99
    neuron_patterns[100] = 16'h170A;  // Neuron 100
    neuron_patterns[101] = 16'h8010;  // Neuron 101
    neuron_patterns[102] = 16'h4860;  // Neuron 102
    neuron_patterns[103] = 16'h30B4;  // Neuron 103
    neuron_patterns[104] = 16'h4A40;  // Neuron 104
    neuron_patterns[105] = 16'h591C;  // Neuron 105
    neuron_patterns[106] = 16'hBC28;  // Neuron 106
    neuron_patterns[107] = 16'h0F48;  // Neuron 107
    neuron_patterns[108] = 16'hE624;  // Neuron 108
    neuron_patterns[109] = 16'h66B3;  // Neuron 109
    neuron_patterns[110] = 16'h242C;  // Neuron 110
    neuron_patterns[111] = 16'h0208;  // Neuron 111
    neuron_patterns[112] = 16'h0C30;  // Neuron 112
    neuron_patterns[113] = 16'hB000;  // Neuron 113
    neuron_patterns[114] = 16'h2022;  // Neuron 114
    neuron_patterns[115] = 16'hA252;  // Neuron 115
    neuron_patterns[116] = 16'h9421;  // Neuron 116
    neuron_patterns[117] = 16'h8210;  // Neuron 117
    neuron_patterns[118] = 16'h2418;  // Neuron 118
    neuron_patterns[119] = 16'h1115;  // Neuron 119
    neuron_patterns[120] = 16'h0101;  // Neuron 120
    neuron_patterns[121] = 16'h4500;  // Neuron 121
    neuron_patterns[122] = 16'h21C0;  // Neuron 122
    neuron_patterns[123] = 16'h3B28;  // Neuron 123
    neuron_patterns[124] = 16'h930A;  // Neuron 124
    neuron_patterns[125] = 16'h0010;  // Neuron 125
    neuron_patterns[126] = 16'h0861;  // Neuron 126
    neuron_patterns[127] = 16'h3060;  // Neuron 127
    neuron_patterns[128] = 16'h4A00;  // Neuron 128
    neuron_patterns[129] = 16'hC008;  // Neuron 129
    neuron_patterns[130] = 16'h35A8;  // Neuron 130
    neuron_patterns[131] = 16'h0B40;  // Neuron 131
    neuron_patterns[132] = 16'hE300;  // Neuron 132
    neuron_patterns[133] = 16'h2003;  // Neuron 133
    neuron_patterns[134] = 16'h3020;  // Neuron 134
    neuron_patterns[135] = 16'h6681;  // Neuron 135
    neuron_patterns[136] = 16'h8C40;  // Neuron 136
    neuron_patterns[137] = 16'h8000;  // Neuron 137
    neuron_patterns[138] = 16'hA000;  // Neuron 138
    neuron_patterns[139] = 16'h8858;  // Neuron 139
    neuron_patterns[140] = 16'h9419;  // Neuron 140
    neuron_patterns[141] = 16'h9512;  // Neuron 141
    neuron_patterns[142] = 16'h0108;  // Neuron 142
    neuron_patterns[143] = 16'h5101;  // Neuron 143
    neuron_patterns[144] = 16'h0201;  // Neuron 144
    neuron_patterns[145] = 16'h6580;  // Neuron 145
    neuron_patterns[146] = 16'h0240;  // Neuron 146
    neuron_patterns[147] = 16'hCD00;  // Neuron 147
    neuron_patterns[148] = 16'h1002;  // Neuron 148
    neuron_patterns[149] = 16'h0010;  // Neuron 149
    neuron_patterns[150] = 16'h0040;  // Neuron 150
    neuron_patterns[151] = 16'h0000;  // Neuron 151
    neuron_patterns[152] = 16'h42C2;  // Neuron 152
    neuron_patterns[153] = 16'h5988;  // Neuron 153
    neuron_patterns[154] = 16'h3828;  // Neuron 154
    neuron_patterns[155] = 16'h0A40;  // Neuron 155
    neuron_patterns[156] = 16'hA214;  // Neuron 156
    neuron_patterns[157] = 16'h2233;  // Neuron 157
    neuron_patterns[158] = 16'hA02C;  // Neuron 158
    neuron_patterns[159] = 16'h0201;  // Neuron 159
    neuron_patterns[160] = 16'h0C28;  // Neuron 160
    neuron_patterns[161] = 16'h9000;  // Neuron 161
    neuron_patterns[162] = 16'hA812;  // Neuron 162
    neuron_patterns[163] = 16'h8052;  // Neuron 163
    neuron_patterns[164] = 16'h9018;  // Neuron 164
    neuron_patterns[165] = 16'h0202;  // Neuron 165
    neuron_patterns[166] = 16'h2400;  // Neuron 166
    neuron_patterns[167] = 16'h4201;  // Neuron 167
    neuron_patterns[168] = 16'h0001;  // Neuron 168
    neuron_patterns[169] = 16'h6D84;  // Neuron 169
    neuron_patterns[170] = 16'h0A40;  // Neuron 170
    neuron_patterns[171] = 16'h8730;  // Neuron 171
    neuron_patterns[172] = 16'h1422;  // Neuron 172
    neuron_patterns[173] = 16'h8010;  // Neuron 173
    neuron_patterns[174] = 16'h0255;  // Neuron 174
    neuron_patterns[175] = 16'h3180;  // Neuron 175
    neuron_patterns[176] = 16'h4E80;  // Neuron 176
    neuron_patterns[177] = 16'h711D;  // Neuron 177
    neuron_patterns[178] = 16'h2C29;  // Neuron 178
    neuron_patterns[179] = 16'h8D41;  // Neuron 179
    neuron_patterns[180] = 16'h8310;  // Neuron 180
    neuron_patterns[181] = 16'h6433;  // Neuron 181
    neuron_patterns[182] = 16'hA028;  // Neuron 182
    neuron_patterns[183] = 16'h0F05;  // Neuron 183
    neuron_patterns[184] = 16'h0020;  // Neuron 184
    neuron_patterns[185] = 16'h8000;  // Neuron 185
    neuron_patterns[186] = 16'hAC02;  // Neuron 186
    neuron_patterns[187] = 16'h8092;  // Neuron 187
    neuron_patterns[188] = 16'h9412;  // Neuron 188
    neuron_patterns[189] = 16'hAA22;  // Neuron 189
    neuron_patterns[190] = 16'h0648;  // Neuron 190
    neuron_patterns[191] = 16'h4B57;  // Neuron 191
    neuron_patterns[192] = 16'h4203;  // Neuron 192
    neuron_patterns[193] = 16'h4500;  // Neuron 193
    neuron_patterns[194] = 16'h0B60;  // Neuron 194
    neuron_patterns[195] = 16'h9BB8;  // Neuron 195
    neuron_patterns[196] = 16'h970A;  // Neuron 196
    neuron_patterns[197] = 16'h9014;  // Neuron 197
    neuron_patterns[198] = 16'h0645;  // Neuron 198
    neuron_patterns[199] = 16'h118C;  // Neuron 199
    neuron_patterns[200] = 16'h5E11;  // Neuron 200
    neuron_patterns[201] = 16'hF91F;  // Neuron 201
    neuron_patterns[202] = 16'hBC29;  // Neuron 202
    neuron_patterns[203] = 16'h0B41;  // Neuron 203
    neuron_patterns[204] = 16'hA294;  // Neuron 204
    neuron_patterns[205] = 16'h7037;  // Neuron 205
    neuron_patterns[206] = 16'hE028;  // Neuron 206
    neuron_patterns[207] = 16'h6320;  // Neuron 207
    neuron_patterns[208] = 16'h2C30;  // Neuron 208
    neuron_patterns[209] = 16'h8000;  // Neuron 209
    neuron_patterns[210] = 16'hACB2;  // Neuron 210
    neuron_patterns[211] = 16'h8052;  // Neuron 211
    neuron_patterns[212] = 16'h9031;  // Neuron 212
    neuron_patterns[213] = 16'h8602;  // Neuron 213
    neuron_patterns[214] = 16'h4450;  // Neuron 214
    neuron_patterns[215] = 16'hCB51;  // Neuron 215
    neuron_patterns[216] = 16'h0121;  // Neuron 216
    neuron_patterns[217] = 16'h4500;  // Neuron 217
    neuron_patterns[218] = 16'h0940;  // Neuron 218
    neuron_patterns[219] = 16'h93C8;  // Neuron 219
    neuron_patterns[220] = 16'h8212;  // Neuron 220
    neuron_patterns[221] = 16'h9034;  // Neuron 221
    neuron_patterns[222] = 16'h0044;  // Neuron 222
    neuron_patterns[223] = 16'h30CC;  // Neuron 223
    neuron_patterns[224] = 16'h4620;  // Neuron 224
    neuron_patterns[225] = 16'hF11D;  // Neuron 225
    neuron_patterns[226] = 16'hBC01;  // Neuron 226
    neuron_patterns[227] = 16'h0B40;  // Neuron 227
    neuron_patterns[228] = 16'hA284;  // Neuron 228
    neuron_patterns[229] = 16'h7211;  // Neuron 229
    neuron_patterns[230] = 16'h0008;  // Neuron 230
    neuron_patterns[231] = 16'h2228;  // Neuron 231
    neuron_patterns[232] = 16'h0020;  // Neuron 232
    neuron_patterns[233] = 16'h0000;  // Neuron 233
    neuron_patterns[234] = 16'hB432;  // Neuron 234
    neuron_patterns[235] = 16'h80D0;  // Neuron 235
    neuron_patterns[236] = 16'h9014;  // Neuron 236
    neuron_patterns[237] = 16'h8622;  // Neuron 237
    neuron_patterns[238] = 16'h4408;  // Neuron 238
    neuron_patterns[239] = 16'hCB53;  // Neuron 239
    neuron_patterns[240] = 16'h0B21;  // Neuron 240
    neuron_patterns[241] = 16'h4504;  // Neuron 241
    neuron_patterns[242] = 16'h8140;  // Neuron 242
    neuron_patterns[243] = 16'h93C8;  // Neuron 243
    neuron_patterns[244] = 16'h924A;  // Neuron 244
    neuron_patterns[245] = 16'h0004;  // Neuron 245
    neuron_patterns[246] = 16'h0040;  // Neuron 246
    neuron_patterns[247] = 16'h3084;  // Neuron 247
    neuron_patterns[248] = 16'h4A00;  // Neuron 248
    neuron_patterns[249] = 16'h7008;  // Neuron 249
    neuron_patterns[250] = 16'hBCA8;  // Neuron 250
    neuron_patterns[251] = 16'h0B60;  // Neuron 251
    neuron_patterns[252] = 16'hE300;  // Neuron 252
    neuron_patterns[253] = 16'h6233;  // Neuron 253
    neuron_patterns[254] = 16'h0004;  // Neuron 254
    neuron_patterns[255] = 16'h2200;  // Neuron 255
  end

endmodule
