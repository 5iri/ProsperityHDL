// ProsperityHDL Tile Data (256x16)
// Generated from SDT CIFAR-10 data
module fc_q_enc_1_tile_data;

  // Tile memory: 256 rows x 16 bits
  reg [15:0] tile_memory [0:255];

  initial begin
    tile_memory[  0] = 16'h04E0;
    tile_memory[  1] = 16'h69F8;
    tile_memory[  2] = 16'h5EFA;
    tile_memory[  3] = 16'hE22B;
    tile_memory[  4] = 16'h8E97;
    tile_memory[  5] = 16'h86B9;
    tile_memory[  6] = 16'hC211;
    tile_memory[  7] = 16'hF0AC;
    tile_memory[  8] = 16'h3950;
    tile_memory[  9] = 16'hD931;
    tile_memory[ 10] = 16'h4077;
    tile_memory[ 11] = 16'hF92B;
    tile_memory[ 12] = 16'h3AC2;
    tile_memory[ 13] = 16'hDB04;
    tile_memory[ 14] = 16'h6FD2;
    tile_memory[ 15] = 16'h90E4;
    tile_memory[ 16] = 16'hFF13;
    tile_memory[ 17] = 16'h0135;
    tile_memory[ 18] = 16'hE294;
    tile_memory[ 19] = 16'h66F3;
    tile_memory[ 20] = 16'h1A60;
    tile_memory[ 21] = 16'hF596;
    tile_memory[ 22] = 16'h0702;
    tile_memory[ 23] = 16'h3E0D;
    tile_memory[ 24] = 16'h4851;
    tile_memory[ 25] = 16'h8941;
    tile_memory[ 26] = 16'h1C01;
    tile_memory[ 27] = 16'h09CB;
    tile_memory[ 28] = 16'h44BB;
    tile_memory[ 29] = 16'h3EA2;
    tile_memory[ 30] = 16'h9DC9;
    tile_memory[ 31] = 16'hA12D;
    tile_memory[ 32] = 16'h40AA;
    tile_memory[ 33] = 16'hD4F9;
    tile_memory[ 34] = 16'h0154;
    tile_memory[ 35] = 16'hD00F;
    tile_memory[ 36] = 16'h41E0;
    tile_memory[ 37] = 16'h870D;
    tile_memory[ 38] = 16'h6342;
    tile_memory[ 39] = 16'h61B0;
    tile_memory[ 40] = 16'h30C3;
    tile_memory[ 41] = 16'hDA9C;
    tile_memory[ 42] = 16'hEB93;
    tile_memory[ 43] = 16'hCC01;
    tile_memory[ 44] = 16'hD940;
    tile_memory[ 45] = 16'hBB94;
    tile_memory[ 46] = 16'hCB77;
    tile_memory[ 47] = 16'h9EDB;
    tile_memory[ 48] = 16'h9086;
    tile_memory[ 49] = 16'h6046;
    tile_memory[ 50] = 16'h9725;
    tile_memory[ 51] = 16'h6DB0;
    tile_memory[ 52] = 16'hE16D;
    tile_memory[ 53] = 16'h5032;
    tile_memory[ 54] = 16'hB627;
    tile_memory[ 55] = 16'h1D46;
    tile_memory[ 56] = 16'hC684;
    tile_memory[ 57] = 16'h74EB;
    tile_memory[ 58] = 16'hE617;
    tile_memory[ 59] = 16'h7B99;
    tile_memory[ 60] = 16'hD12F;
    tile_memory[ 61] = 16'h2832;
    tile_memory[ 62] = 16'hA66E;
    tile_memory[ 63] = 16'hB2DD;
    tile_memory[ 64] = 16'h1C31;
    tile_memory[ 65] = 16'hA5B8;
    tile_memory[ 66] = 16'h78AC;
    tile_memory[ 67] = 16'h1CBC;
    tile_memory[ 68] = 16'h0280;
    tile_memory[ 69] = 16'h28A4;
    tile_memory[ 70] = 16'h540F;
    tile_memory[ 71] = 16'h91AB;
    tile_memory[ 72] = 16'hA835;
    tile_memory[ 73] = 16'hA94E;
    tile_memory[ 74] = 16'hF002;
    tile_memory[ 75] = 16'hA0EE;
    tile_memory[ 76] = 16'hB679;
    tile_memory[ 77] = 16'h18DA;
    tile_memory[ 78] = 16'h0B92;
    tile_memory[ 79] = 16'h1FC8;
    tile_memory[ 80] = 16'hAFCB;
    tile_memory[ 81] = 16'hF417;
    tile_memory[ 82] = 16'h9C5D;
    tile_memory[ 83] = 16'h5018;
    tile_memory[ 84] = 16'hEACD;
    tile_memory[ 85] = 16'h0F4E;
    tile_memory[ 86] = 16'hC44A;
    tile_memory[ 87] = 16'h9D9F;
    tile_memory[ 88] = 16'hFA1D;
    tile_memory[ 89] = 16'hD65E;
    tile_memory[ 90] = 16'h08C8;
    tile_memory[ 91] = 16'hA468;
    tile_memory[ 92] = 16'h98D9;
    tile_memory[ 93] = 16'h72C9;
    tile_memory[ 94] = 16'h9582;
    tile_memory[ 95] = 16'hE9D3;
    tile_memory[ 96] = 16'h88D0;
    tile_memory[ 97] = 16'h0582;
    tile_memory[ 98] = 16'h3B72;
    tile_memory[ 99] = 16'hEA9E;
    tile_memory[100] = 16'h151D;
    tile_memory[101] = 16'h617E;
    tile_memory[102] = 16'h0623;
    tile_memory[103] = 16'h312C;
    tile_memory[104] = 16'h46AA;
    tile_memory[105] = 16'hC725;
    tile_memory[106] = 16'h83B4;
    tile_memory[107] = 16'h19E2;
    tile_memory[108] = 16'h7320;
    tile_memory[109] = 16'h31B4;
    tile_memory[110] = 16'h9390;
    tile_memory[111] = 16'h6FDE;
    tile_memory[112] = 16'h8B74;
    tile_memory[113] = 16'h7264;
    tile_memory[114] = 16'h0381;
    tile_memory[115] = 16'h8625;
    tile_memory[116] = 16'hDE23;
    tile_memory[117] = 16'h0F79;
    tile_memory[118] = 16'h6EB4;
    tile_memory[119] = 16'h235D;
    tile_memory[120] = 16'hE1E6;
    tile_memory[121] = 16'hE8C0;
    tile_memory[122] = 16'hB415;
    tile_memory[123] = 16'hA966;
    tile_memory[124] = 16'h78E4;
    tile_memory[125] = 16'h764E;
    tile_memory[126] = 16'hD216;
    tile_memory[127] = 16'hAF64;
    tile_memory[128] = 16'h9657;
    tile_memory[129] = 16'h0B31;
    tile_memory[130] = 16'hB200;
    tile_memory[131] = 16'hB08E;
    tile_memory[132] = 16'h86AE;
    tile_memory[133] = 16'hAE25;
    tile_memory[134] = 16'h3196;
    tile_memory[135] = 16'h1735;
    tile_memory[136] = 16'h546C;
    tile_memory[137] = 16'h1C4A;
    tile_memory[138] = 16'h88E3;
    tile_memory[139] = 16'h3C73;
    tile_memory[140] = 16'h406C;
    tile_memory[141] = 16'h7C57;
    tile_memory[142] = 16'h8894;
    tile_memory[143] = 16'h8B19;
    tile_memory[144] = 16'hC45A;
    tile_memory[145] = 16'hCACD;
    tile_memory[146] = 16'hF0EE;
    tile_memory[147] = 16'hE466;
    tile_memory[148] = 16'hEA3A;
    tile_memory[149] = 16'h3EF1;
    tile_memory[150] = 16'h1565;
    tile_memory[151] = 16'h74E6;
    tile_memory[152] = 16'hDA4F;
    tile_memory[153] = 16'hF58A;
    tile_memory[154] = 16'hDAF8;
    tile_memory[155] = 16'h5BF0;
    tile_memory[156] = 16'h3BE5;
    tile_memory[157] = 16'h174E;
    tile_memory[158] = 16'hEC17;
    tile_memory[159] = 16'h7FF7;
    tile_memory[160] = 16'h1E42;
    tile_memory[161] = 16'h17F9;
    tile_memory[162] = 16'hF4DF;
    tile_memory[163] = 16'h8ABE;
    tile_memory[164] = 16'h79FF;
    tile_memory[165] = 16'hEC79;
    tile_memory[166] = 16'h3723;
    tile_memory[167] = 16'hD09B;
    tile_memory[168] = 16'h84BB;
    tile_memory[169] = 16'hDD6E;
    tile_memory[170] = 16'h1DAB;
    tile_memory[171] = 16'hE4C7;
    tile_memory[172] = 16'hB46B;
    tile_memory[173] = 16'h94D4;
    tile_memory[174] = 16'h98D3;
    tile_memory[175] = 16'h4811;
    tile_memory[176] = 16'hA01D;
    tile_memory[177] = 16'h9A5D;
    tile_memory[178] = 16'h5AF2;
    tile_memory[179] = 16'hFF8D;
    tile_memory[180] = 16'hC3BE;
    tile_memory[181] = 16'h2CF8;
    tile_memory[182] = 16'h9167;
    tile_memory[183] = 16'hFBD8;
    tile_memory[184] = 16'h6B34;
    tile_memory[185] = 16'h5DEE;
    tile_memory[186] = 16'hBE4F;
    tile_memory[187] = 16'hCD67;
    tile_memory[188] = 16'h1C49;
    tile_memory[189] = 16'hD0E8;
    tile_memory[190] = 16'h6CB3;
    tile_memory[191] = 16'hFB0F;
    tile_memory[192] = 16'h9E5F;
    tile_memory[193] = 16'h77F2;
    tile_memory[194] = 16'h85FB;
    tile_memory[195] = 16'hE8D7;
    tile_memory[196] = 16'h4FDF;
    tile_memory[197] = 16'h8FBF;
    tile_memory[198] = 16'hCDED;
    tile_memory[199] = 16'hCFAB;
    tile_memory[200] = 16'hB3D7;
    tile_memory[201] = 16'hD31F;
    tile_memory[202] = 16'h9A6A;
    tile_memory[203] = 16'h3CF7;
    tile_memory[204] = 16'hAE2D;
    tile_memory[205] = 16'hB5B0;
    tile_memory[206] = 16'h6914;
    tile_memory[207] = 16'hCEA8;
    tile_memory[208] = 16'hE2C2;
    tile_memory[209] = 16'hBBEF;
    tile_memory[210] = 16'hFD77;
    tile_memory[211] = 16'h7365;
    tile_memory[212] = 16'h577E;
    tile_memory[213] = 16'hFDB1;
    tile_memory[214] = 16'hEE73;
    tile_memory[215] = 16'h4CDF;
    tile_memory[216] = 16'h7883;
    tile_memory[217] = 16'hFDFD;
    tile_memory[218] = 16'hEAC9;
    tile_memory[219] = 16'h6573;
    tile_memory[220] = 16'h9EF3;
    tile_memory[221] = 16'hDB7A;
    tile_memory[222] = 16'h621E;
    tile_memory[223] = 16'h843D;
    tile_memory[224] = 16'h627F;
    tile_memory[225] = 16'h4DC1;
    tile_memory[226] = 16'hD0CA;
    tile_memory[227] = 16'h6C7F;
    tile_memory[228] = 16'h7BFD;
    tile_memory[229] = 16'hF4CC;
    tile_memory[230] = 16'h95DD;
    tile_memory[231] = 16'h4E70;
    tile_memory[232] = 16'hCB4C;
    tile_memory[233] = 16'h6F71;
    tile_memory[234] = 16'h722E;
    tile_memory[235] = 16'h502F;
    tile_memory[236] = 16'h22FC;
    tile_memory[237] = 16'hBF65;
    tile_memory[238] = 16'h0917;
    tile_memory[239] = 16'h863E;
    tile_memory[240] = 16'hD6D8;
    tile_memory[241] = 16'h41B5;
    tile_memory[242] = 16'h751C;
    tile_memory[243] = 16'h1495;
    tile_memory[244] = 16'h2F75;
    tile_memory[245] = 16'hF370;
    tile_memory[246] = 16'h53E8;
    tile_memory[247] = 16'h94DF;
    tile_memory[248] = 16'hD603;
    tile_memory[249] = 16'hFEE6;
    tile_memory[250] = 16'h2866;
    tile_memory[251] = 16'h0F86;
    tile_memory[252] = 16'h7179;
    tile_memory[253] = 16'h465A;
    tile_memory[254] = 16'hF71F;
    tile_memory[255] = 16'h0CE4;
  end

endmodule
