// ProSparsity Hardware Test Data
// Raw spike patterns: 256 neurons × 16 timesteps
module fc_k_enc_7_tile_data;

  // Neuron spike patterns: 256 neurons × 16 timesteps
  reg [15:0] neuron_patterns [0:255];

  initial begin
    neuron_patterns[  0] = 16'h5AA0;  // Neuron 0
    neuron_patterns[  1] = 16'h69FE;  // Neuron 1
    neuron_patterns[  2] = 16'hDFFF;  // Neuron 2
    neuron_patterns[  3] = 16'hFB79;  // Neuron 3
    neuron_patterns[  4] = 16'h8FFF;  // Neuron 4
    neuron_patterns[  5] = 16'hFBB9;  // Neuron 5
    neuron_patterns[  6] = 16'hDAD9;  // Neuron 6
    neuron_patterns[  7] = 16'hFFB7;  // Neuron 7
    neuron_patterns[  8] = 16'hE971;  // Neuron 8
    neuron_patterns[  9] = 16'hDBF5;  // Neuron 9
    neuron_patterns[ 10] = 16'h48F7;  // Neuron 10
    neuron_patterns[ 11] = 16'hCFBB;  // Neuron 11
    neuron_patterns[ 12] = 16'h3FF7;  // Neuron 12
    neuron_patterns[ 13] = 16'hDF4C;  // Neuron 13
    neuron_patterns[ 14] = 16'h6FD3;  // Neuron 14
    neuron_patterns[ 15] = 16'hF6E0;  // Neuron 15
    neuron_patterns[ 16] = 16'hFF1A;  // Neuron 16
    neuron_patterns[ 17] = 16'h2335;  // Neuron 17
    neuron_patterns[ 18] = 16'hF296;  // Neuron 18
    neuron_patterns[ 19] = 16'hF6F3;  // Neuron 19
    neuron_patterns[ 20] = 16'h1EAB;  // Neuron 20
    neuron_patterns[ 21] = 16'hD7DE;  // Neuron 21
    neuron_patterns[ 22] = 16'h7F06;  // Neuron 22
    neuron_patterns[ 23] = 16'hFE7D;  // Neuron 23
    neuron_patterns[ 24] = 16'hCD5D;  // Neuron 24
    neuron_patterns[ 25] = 16'hDF42;  // Neuron 25
    neuron_patterns[ 26] = 16'h3D13;  // Neuron 26
    neuron_patterns[ 27] = 16'h0BFB;  // Neuron 27
    neuron_patterns[ 28] = 16'h5DDF;  // Neuron 28
    neuron_patterns[ 29] = 16'hB7AF;  // Neuron 29
    neuron_patterns[ 30] = 16'hBD4D;  // Neuron 30
    neuron_patterns[ 31] = 16'h613F;  // Neuron 31
    neuron_patterns[ 32] = 16'h62FA;  // Neuron 32
    neuron_patterns[ 33] = 16'hDCF9;  // Neuron 33
    neuron_patterns[ 34] = 16'h8955;  // Neuron 34
    neuron_patterns[ 35] = 16'hDE2F;  // Neuron 35
    neuron_patterns[ 36] = 16'h71F8;  // Neuron 36
    neuron_patterns[ 37] = 16'hA7AC;  // Neuron 37
    neuron_patterns[ 38] = 16'h67E7;  // Neuron 38
    neuron_patterns[ 39] = 16'hE76D;  // Neuron 39
    neuron_patterns[ 40] = 16'hBFD3;  // Neuron 40
    neuron_patterns[ 41] = 16'hDAB9;  // Neuron 41
    neuron_patterns[ 42] = 16'hEB8B;  // Neuron 42
    neuron_patterns[ 43] = 16'hDD29;  // Neuron 43
    neuron_patterns[ 44] = 16'hF9F0;  // Neuron 44
    neuron_patterns[ 45] = 16'h939C;  // Neuron 45
    neuron_patterns[ 46] = 16'h7F77;  // Neuron 46
    neuron_patterns[ 47] = 16'hAEBF;  // Neuron 47
    neuron_patterns[ 48] = 16'h5AF4;  // Neuron 48
    neuron_patterns[ 49] = 16'hF7E6;  // Neuron 49
    neuron_patterns[ 50] = 16'hFD77;  // Neuron 50
    neuron_patterns[ 51] = 16'h7B5A;  // Neuron 51
    neuron_patterns[ 52] = 16'h976E;  // Neuron 52
    neuron_patterns[ 53] = 16'hFBF1;  // Neuron 53
    neuron_patterns[ 54] = 16'hDBCB;  // Neuron 54
    neuron_patterns[ 55] = 16'hFF8B;  // Neuron 55
    neuron_patterns[ 56] = 16'hC9CB;  // Neuron 56
    neuron_patterns[ 57] = 16'hC7E5;  // Neuron 57
    neuron_patterns[ 58] = 16'h2DD6;  // Neuron 58
    neuron_patterns[ 59] = 16'h6713;  // Neuron 59
    neuron_patterns[ 60] = 16'hAFBB;  // Neuron 60
    neuron_patterns[ 61] = 16'h97CC;  // Neuron 61
    neuron_patterns[ 62] = 16'hA859;  // Neuron 62
    neuron_patterns[ 63] = 16'hE566;  // Neuron 63
    neuron_patterns[ 64] = 16'hE71C;  // Neuron 64
    neuron_patterns[ 65] = 16'h4653;  // Neuron 65
    neuron_patterns[ 66] = 16'hF9C3;  // Neuron 66
    neuron_patterns[ 67] = 16'hD462;  // Neuron 67
    neuron_patterns[ 68] = 16'h2FAA;  // Neuron 68
    neuron_patterns[ 69] = 16'hDBDC;  // Neuron 69
    neuron_patterns[ 70] = 16'h7F0E;  // Neuron 70
    neuron_patterns[ 71] = 16'hD4F3;  // Neuron 71
    neuron_patterns[ 72] = 16'hDFAC;  // Neuron 72
    neuron_patterns[ 73] = 16'hD713;  // Neuron 73
    neuron_patterns[ 74] = 16'h7F12;  // Neuron 74
    neuron_patterns[ 75] = 16'h33FF;  // Neuron 75
    neuron_patterns[ 76] = 16'hD9CF;  // Neuron 76
    neuron_patterns[ 77] = 16'hA93B;  // Neuron 77
    neuron_patterns[ 78] = 16'hBF7E;  // Neuron 78
    neuron_patterns[ 79] = 16'hE8AF;  // Neuron 79
    neuron_patterns[ 80] = 16'h6FB2;  // Neuron 80
    neuron_patterns[ 81] = 16'hEFF8;  // Neuron 81
    neuron_patterns[ 82] = 16'hECD7;  // Neuron 82
    neuron_patterns[ 83] = 16'hCF15;  // Neuron 83
    neuron_patterns[ 84] = 16'h70B0;  // Neuron 84
    neuron_patterns[ 85] = 16'hF3B8;  // Neuron 85
    neuron_patterns[ 86] = 16'hADEF;  // Neuron 86
    neuron_patterns[ 87] = 16'hEF1D;  // Neuron 87
    neuron_patterns[ 88] = 16'hAFAF;  // Neuron 88
    neuron_patterns[ 89] = 16'h9BAB;  // Neuron 89
    neuron_patterns[ 90] = 16'hB38F;  // Neuron 90
    neuron_patterns[ 91] = 16'h7B3F;  // Neuron 91
    neuron_patterns[ 92] = 16'hD9B8;  // Neuron 92
    neuron_patterns[ 93] = 16'hEEBD;  // Neuron 93
    neuron_patterns[ 94] = 16'h7E3B;  // Neuron 94
    neuron_patterns[ 95] = 16'hEEBF;  // Neuron 95
    neuron_patterns[ 96] = 16'hFAC2;  // Neuron 96
    neuron_patterns[ 97] = 16'h5BFE;  // Neuron 97
    neuron_patterns[ 98] = 16'hDF19;  // Neuron 98
    neuron_patterns[ 99] = 16'hFFFF;  // Neuron 99
    neuron_patterns[100] = 16'hBD6F;  // Neuron 100
    neuron_patterns[101] = 16'hFBB7;  // Neuron 101
    neuron_patterns[102] = 16'hFADB;  // Neuron 102
    neuron_patterns[103] = 16'hD74B;  // Neuron 103
    neuron_patterns[104] = 16'hEBF9;  // Neuron 104
    neuron_patterns[105] = 16'hD3AF;  // Neuron 105
    neuron_patterns[106] = 16'hF8F3;  // Neuron 106
    neuron_patterns[107] = 16'h8F3B;  // Neuron 107
    neuron_patterns[108] = 16'h7F3F;  // Neuron 108
    neuron_patterns[109] = 16'hA68E;  // Neuron 109
    neuron_patterns[110] = 16'hED15;  // Neuron 110
    neuron_patterns[111] = 16'hF6F9;  // Neuron 111
    neuron_patterns[112] = 16'h579D;  // Neuron 112
    neuron_patterns[113] = 16'h64F3;  // Neuron 113
    neuron_patterns[114] = 16'h3BF2;  // Neuron 114
    neuron_patterns[115] = 16'hF776;  // Neuron 115
    neuron_patterns[116] = 16'h0DFB;  // Neuron 116
    neuron_patterns[117] = 16'hC6FC;  // Neuron 117
    neuron_patterns[118] = 16'hFEB6;  // Neuron 118
    neuron_patterns[119] = 16'hF17E;  // Neuron 119
    neuron_patterns[120] = 16'hE776;  // Neuron 120
    neuron_patterns[121] = 16'hDF57;  // Neuron 121
    neuron_patterns[122] = 16'hED10;  // Neuron 122
    neuron_patterns[123] = 16'h3AF1;  // Neuron 123
    neuron_patterns[124] = 16'hDBFD;  // Neuron 124
    neuron_patterns[125] = 16'hEBE7;  // Neuron 125
    neuron_patterns[126] = 16'hBFED;  // Neuron 126
    neuron_patterns[127] = 16'hC77F;  // Neuron 127
    neuron_patterns[128] = 16'hFFDE;  // Neuron 128
    neuron_patterns[129] = 16'hFEF8;  // Neuron 129
    neuron_patterns[130] = 16'hBA4D;  // Neuron 130
    neuron_patterns[131] = 16'hFF74;  // Neuron 131
    neuron_patterns[132] = 16'h77B3;  // Neuron 132
    neuron_patterns[133] = 16'hABAE;  // Neuron 133
    neuron_patterns[134] = 16'hF5E7;  // Neuron 134
    neuron_patterns[135] = 16'hFFDE;  // Neuron 135
    neuron_patterns[136] = 16'hEFAD;  // Neuron 136
    neuron_patterns[137] = 16'hDCFB;  // Neuron 137
    neuron_patterns[138] = 16'h2FCA;  // Neuron 138
    neuron_patterns[139] = 16'hFB3F;  // Neuron 139
    neuron_patterns[140] = 16'hF9BF;  // Neuron 140
    neuron_patterns[141] = 16'hD2FF;  // Neuron 141
    neuron_patterns[142] = 16'h757C;  // Neuron 142
    neuron_patterns[143] = 16'hAFE7;  // Neuron 143
    neuron_patterns[144] = 16'h7FE0;  // Neuron 144
    neuron_patterns[145] = 16'hFD86;  // Neuron 145
    neuron_patterns[146] = 16'hDF39;  // Neuron 146
    neuron_patterns[147] = 16'h795A;  // Neuron 147
    neuron_patterns[148] = 16'hFDE5;  // Neuron 148
    neuron_patterns[149] = 16'hFBE4;  // Neuron 149
    neuron_patterns[150] = 16'hDFFF;  // Neuron 150
    neuron_patterns[151] = 16'hE7D3;  // Neuron 151
    neuron_patterns[152] = 16'hFF28;  // Neuron 152
    neuron_patterns[153] = 16'hCA3F;  // Neuron 153
    neuron_patterns[154] = 16'hD9CE;  // Neuron 154
    neuron_patterns[155] = 16'h17B3;  // Neuron 155
    neuron_patterns[156] = 16'h3D75;  // Neuron 156
    neuron_patterns[157] = 16'hA44F;  // Neuron 157
    neuron_patterns[158] = 16'h4B79;  // Neuron 158
    neuron_patterns[159] = 16'hE3FB;  // Neuron 159
    neuron_patterns[160] = 16'h3DFD;  // Neuron 160
    neuron_patterns[161] = 16'h21F5;  // Neuron 161
    neuron_patterns[162] = 16'h3196;  // Neuron 162
    neuron_patterns[163] = 16'hDD6A;  // Neuron 163
    neuron_patterns[164] = 16'h6DEA;  // Neuron 164
    neuron_patterns[165] = 16'hF57A;  // Neuron 165
    neuron_patterns[166] = 16'h7C6D;  // Neuron 166
    neuron_patterns[167] = 16'hDBF5;  // Neuron 167
    neuron_patterns[168] = 16'hC7E4;  // Neuron 168
    neuron_patterns[169] = 16'h5EDA;  // Neuron 169
    neuron_patterns[170] = 16'h6F13;  // Neuron 170
    neuron_patterns[171] = 16'hA2EB;  // Neuron 171
    neuron_patterns[172] = 16'h7DFD;  // Neuron 172
    neuron_patterns[173] = 16'hB54B;  // Neuron 173
    neuron_patterns[174] = 16'hBD7E;  // Neuron 174
    neuron_patterns[175] = 16'h7B63;  // Neuron 175
    neuron_patterns[176] = 16'h56D7;  // Neuron 176
    neuron_patterns[177] = 16'h9EFA;  // Neuron 177
    neuron_patterns[178] = 16'hB37F;  // Neuron 178
    neuron_patterns[179] = 16'h7F66;  // Neuron 179
    neuron_patterns[180] = 16'hF938;  // Neuron 180
    neuron_patterns[181] = 16'hF7BA;  // Neuron 181
    neuron_patterns[182] = 16'hFD77;  // Neuron 182
    neuron_patterns[183] = 16'hDB4F;  // Neuron 183
    neuron_patterns[184] = 16'hFF55;  // Neuron 184
    neuron_patterns[185] = 16'h9EE9;  // Neuron 185
    neuron_patterns[186] = 16'hF38B;  // Neuron 186
    neuron_patterns[187] = 16'hDB69;  // Neuron 187
    neuron_patterns[188] = 16'hFDFD;  // Neuron 188
    neuron_patterns[189] = 16'h13DC;  // Neuron 189
    neuron_patterns[190] = 16'h3DD0;  // Neuron 190
    neuron_patterns[191] = 16'h6FAF;  // Neuron 191
    neuron_patterns[192] = 16'hFA8B;  // Neuron 192
    neuron_patterns[193] = 16'hC8DB;  // Neuron 193
    neuron_patterns[194] = 16'h8FDD;  // Neuron 194
    neuron_patterns[195] = 16'hD9F4;  // Neuron 195
    neuron_patterns[196] = 16'hFFEF;  // Neuron 196
    neuron_patterns[197] = 16'h7BFA;  // Neuron 197
    neuron_patterns[198] = 16'hFB5D;  // Neuron 198
    neuron_patterns[199] = 16'h478B;  // Neuron 199
    neuron_patterns[200] = 16'h5B3E;  // Neuron 200
    neuron_patterns[201] = 16'hF2ED;  // Neuron 201
    neuron_patterns[202] = 16'hA9DF;  // Neuron 202
    neuron_patterns[203] = 16'hAF17;  // Neuron 203
    neuron_patterns[204] = 16'h357F;  // Neuron 204
    neuron_patterns[205] = 16'hD6BE;  // Neuron 205
    neuron_patterns[206] = 16'h1AB3;  // Neuron 206
    neuron_patterns[207] = 16'hE8E3;  // Neuron 207
    neuron_patterns[208] = 16'hEF5C;  // Neuron 208
    neuron_patterns[209] = 16'h2C99;  // Neuron 209
    neuron_patterns[210] = 16'hB3EB;  // Neuron 210
    neuron_patterns[211] = 16'hDBEB;  // Neuron 211
    neuron_patterns[212] = 16'hCFBE;  // Neuron 212
    neuron_patterns[213] = 16'hEBFC;  // Neuron 213
    neuron_patterns[214] = 16'h7F3C;  // Neuron 214
    neuron_patterns[215] = 16'hD9F3;  // Neuron 215
    neuron_patterns[216] = 16'hF57D;  // Neuron 216
    neuron_patterns[217] = 16'hB7A7;  // Neuron 217
    neuron_patterns[218] = 16'h79F1;  // Neuron 218
    neuron_patterns[219] = 16'hEBF9;  // Neuron 219
    neuron_patterns[220] = 16'h197D;  // Neuron 220
    neuron_patterns[221] = 16'hF953;  // Neuron 221
    neuron_patterns[222] = 16'hBD5C;  // Neuron 222
    neuron_patterns[223] = 16'h64B7;  // Neuron 223
    neuron_patterns[224] = 16'h4EF2;  // Neuron 224
    neuron_patterns[225] = 16'hEBFF;  // Neuron 225
    neuron_patterns[226] = 16'h95EB;  // Neuron 226
    neuron_patterns[227] = 16'h2E6F;  // Neuron 227
    neuron_patterns[228] = 16'h7D77;  // Neuron 228
    neuron_patterns[229] = 16'hFBFB;  // Neuron 229
    neuron_patterns[230] = 16'hF5E5;  // Neuron 230
    neuron_patterns[231] = 16'hE75C;  // Neuron 231
    neuron_patterns[232] = 16'hEFF1;  // Neuron 232
    neuron_patterns[233] = 16'hB8BD;  // Neuron 233
    neuron_patterns[234] = 16'hE7EB;  // Neuron 234
    neuron_patterns[235] = 16'h57BF;  // Neuron 235
    neuron_patterns[236] = 16'hBEB8;  // Neuron 236
    neuron_patterns[237] = 16'h1AFC;  // Neuron 237
    neuron_patterns[238] = 16'h7DC1;  // Neuron 238
    neuron_patterns[239] = 16'hEE57;  // Neuron 239
    neuron_patterns[240] = 16'h5AC0;  // Neuron 240
    neuron_patterns[241] = 16'h41CE;  // Neuron 241
    neuron_patterns[242] = 16'hDF3D;  // Neuron 242
    neuron_patterns[243] = 16'hDF5E;  // Neuron 243
    neuron_patterns[244] = 16'hB564;  // Neuron 244
    neuron_patterns[245] = 16'h7BFB;  // Neuron 245
    neuron_patterns[246] = 16'hFACB;  // Neuron 246
    neuron_patterns[247] = 16'h4713;  // Neuron 247
    neuron_patterns[248] = 16'hE5A7;  // Neuron 248
    neuron_patterns[249] = 16'hFBA7;  // Neuron 249
    neuron_patterns[250] = 16'h28D5;  // Neuron 250
    neuron_patterns[251] = 16'h4F1B;  // Neuron 251
    neuron_patterns[252] = 16'h3DB7;  // Neuron 252
    neuron_patterns[253] = 16'hBC9D;  // Neuron 253
    neuron_patterns[254] = 16'hCC9D;  // Neuron 254
    neuron_patterns[255] = 16'hF761;  // Neuron 255
  end

endmodule
